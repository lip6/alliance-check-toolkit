.model sky130_fd_pr__nfet_01v8__model.0 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.5160869
+ k1 = 0.54086565
+ k2 = -0.026708291
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.1052686
+ nfactor = 2.68453
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0314621
+ ua = -7.5795907e-10
+ ub = 1.57049e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.369451
+ ags = 0.380025
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.1 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.5160869
+ k1 = 0.54086565
+ k2 = -0.026708291
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.1052686
+ nfactor = 2.68453
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0314621
+ ua = -7.5795907e-10
+ ub = 1.57049e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.369451
+ ags = 0.380025
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.2 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.166909460e-01 lvth0 = -4.838883101e-09 wvth0 = -6.033932022e-08 pvth0 = 4.833653817e-13
+ k1 = 5.415453773e-01 lk1 = -5.445149777e-09 wk1 = -6.789927122e-08 pk1 = 5.439265313e-13
+ k2 = -2.711805592e-02 lk2 = 3.282539101e-09 wk2 = 4.093220973e-08 pk2 = -3.278991727e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.049996442e-01 lvoff = -2.154547359e-09 wvoff = -2.686651451e-08 pvoff = 2.152218983e-13
+ nfactor = 2.686034709e+00 lnfactor = -1.205390299e-08 wnfactor = -1.503083041e-07 pnfactor = 1.204087658e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.142325993e-02 lu0 = 3.111395108e-10 wu0 = 3.879809903e-09 pu0 = -3.108032685e-14
+ ua = -7.575504764e-10 lua = -3.273155509e-18 wua = -4.081519935e-17 pua = 3.269618276e-22
+ ub = 1.564807772e-18 lub = 4.551910922e-26 wub = 5.676086919e-25 pub = -4.546991763e-30
+ uc = 4.877037585e-11 luc = 3.778080112e-18 wuc = 4.711144720e-17 puc = -3.773997217e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.361739852e+00 la0 = 6.177235391e-08 wa0 = 7.702814400e-07 pa0 = -6.170559776e-12
+ ags = 3.816712633e-01 lags = -1.318786275e-08 wags = -1.644484186e-07 pags = 1.317361089e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.950752899e-24 lb1 = 1.254404981e-30 wb1 = 1.564202776e-29 pb1 = -1.253049370e-34
+ keta = -8.288371258e-03 lketa = -4.055290119e-09 wketa = -5.056816706e-08 pketa = 4.050907648e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.798002168e-02 lpclm = -3.337615616e-07 wpclm = -4.161899621e-06 ppclm = 3.334008721e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.074731372e-03 lpdiblc2 = -1.019510186e-11 wpdiblc2 = -1.271296502e-10 ppdiblc2 = 1.018408422e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.580421702e+08 lpscbe1 = -2.698040880e+01 wpscbe1 = -3.364370440e+02 ppscbe1 = 2.695125162e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.131867870e-01 lkt1 = 1.255986929e-09 wkt1 = 1.566175415e-08 pkt1 = -1.254629609e-13
+ kt2 = -4.539666594e-02 lkt2 = 6.675302662e-10 wkt2 = 8.323888313e-09 pkt2 = -6.668088796e-14
+ at = 140000.0
+ ute = -1.816357404e+00 lute = 2.369112785e-08 wute = 2.954207655e-07 pute = -2.366552532e-12
+ ua1 = 3.613845672e-10 lua1 = 1.172413201e-16 wua1 = 1.461961658e-15 pua1 = -1.171146198e-20
+ ub1 = -6.204600368e-19 lub1 = -1.534863647e-25 wub1 = -1.913925738e-24 pub1 = 1.533204951e-29
+ uc1 = 1.690921780e-11 luc1 = -8.647681916e-18 wuc1 = -1.078338198e-16 puc1 = 8.638336539e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.3 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.071728966e-01 lvth0 = 3.333597610e-08 wvth0 = 7.402623097e-08 pvth0 = -5.554608993e-14
+ k1 = 5.302997219e-01 lk1 = 3.965876745e-08 wk1 = 1.367515665e-07 pk1 = -2.768841837e-13
+ k2 = -2.048316993e-02 lk2 = -2.332856876e-08 wk2 = -6.801314992e-08 pk2 = 1.090573506e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.376480639e-01 ldsub = 8.964883236e-08 wdsub = 2.232778080e-06 pdsub = -8.955195066e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.094655827e-01 lvoff = 1.575737635e-08 wvoff = 5.573196081e-08 pvoff = -1.160629101e-13
+ nfactor = 2.666085505e+00 lnfactor = 6.795808584e-08 wnfactor = -1.912644030e-07 pnfactor = 1.368353806e-12
+ eta0 = 7.407673693e-02 leta0 = 2.375694058e-08 weta0 = 5.916861913e-07 peta0 = -2.373126692e-12
+ etab = -6.482185296e-02 letab = -2.076843965e-08 wetab = -5.172551119e-07 petab = 2.074599561e-12
+ u0 = 3.194993327e-02 lu0 = -1.801234574e-09 wu0 = 3.764492127e-09 pu0 = -3.061781193e-14
+ ua = -7.771556207e-10 lua = 7.535888247e-17 wua = 1.365337502e-15 pua = -5.312815741e-21
+ ub = 1.668742330e-18 lub = -3.713401575e-25 wub = -2.134683279e-24 pub = 6.291323040e-30
+ uc = 5.890739593e-11 luc = -3.687933810e-17 wuc = -3.280617428e-16 puc = 1.127339656e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.490798641e+00 la0 = -4.558548281e-07 wa0 = -1.699489791e-06 pa0 = 3.735164101e-12
+ ags = 3.647656614e-01 lags = 5.461688862e-08 wags = -7.007562172e-07 pags = 3.468376900e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 4.539228699e-24 lb1 = -9.127417519e-30 wb1 = -3.128405553e-29 pb1 = 6.290554088e-35
+ keta = -1.651832020e-02 lketa = 2.895327386e-08 wketa = 8.733344889e-08 pketa = -1.480031059e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.228164149e-01 lpclm = 2.436875115e-06 wpclm = 8.531224325e-06 ppclm = -1.756931660e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.181986903e-03 lpdiblc2 = -4.403740832e-10 wpdiblc2 = -1.256119770e-08 ppdiblc2 = 5.088879447e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.023678574e+08 lpscbe1 = 1.963173455e+02 wpscbe1 = 6.728740879e+02 ppscbe1 = -1.353005796e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.112536839e-01 lkt1 = -6.497275977e-09 wkt1 = 3.446901913e-08 pkt1 = -2.008948760e-13
+ kt2 = -4.402024159e-02 lkt2 = -4.853013239e-09 wkt2 = -1.654486044e-08 pkt2 = 3.306234138e-14
+ at = 1.381328683e+05 lat = 7.488665797e-03 wat = 1.865113957e-01 pat = -7.480572945e-7
+ ute = -1.757166309e+00 lute = -2.137116870e-07 wute = -1.620152226e-06 pute = 5.316400804e-12
+ ua1 = 6.261329075e-10 lua1 = -9.446076166e-16 wua1 = -5.203440883e-15 pua1 = 1.502204122e-20
+ ub1 = -9.508554259e-19 lub1 = 1.171658836e-24 wub1 = 5.193865106e-24 pub1 = -1.317577850e-29
+ uc1 = -4.824542424e-13 luc1 = 6.110659282e-17 wuc1 = 1.704269561e-16 puc1 = -2.522107706e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.4 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.256581141e-01 lvth0 = -3.833840380e-09 wvth0 = -1.440555601e-07 pvth0 = 3.829697225e-13
+ k1 = 5.525508708e-01 lk1 = -5.083531333e-09 wk1 = -2.534878473e-07 pk1 = 5.078037662e-13
+ k2 = -3.311163166e-02 lk2 = 2.064565301e-09 wk2 = 8.878661258e-08 pk2 = -2.062334167e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.822320387e-01 wdsub = -2.220801299e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.030312872e-01 lvoff = 2.819384981e-09 wvoff = 1.380733451e-07 pvoff = -2.816338128e-13
+ nfactor = 2.691123862e+00 lnfactor = 1.761130745e-08 wnfactor = 1.364137978e-06 pnfactor = -1.759227527e-12
+ eta0 = 8.604364330e-02 leta0 = -3.059472010e-10 weta0 = -6.037112053e-07 peta0 = 3.056165700e-14
+ etab = -7.513627443e-02 letab = -2.834536917e-11 wetab = 5.130723758e-07 petab = 2.831473690e-15
+ u0 = 3.078800555e-02 lu0 = 5.351534303e-10 wu0 = 1.512308431e-08 pu0 = -5.345751007e-14
+ ua = -7.785201420e-10 lua = 7.810264280e-17 wua = 2.603165964e-15 pua = -7.801823884e-21
+ ub = 1.523558700e-18 lub = -7.940694862e-26 wub = -2.950677856e-24 pub = 7.932113512e-30
+ uc = 3.955982554e-11 luc = 2.024485577e-18 wuc = 3.331570204e-16 puc = -2.022297756e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.152059407e+04 lvsat = -3.057589258e-03 wvsat = -1.518950790e-01 pvsat = 3.054284983e-7
+ a0 = 1.249877415e+00 la0 = 2.858620026e-08 wa0 = 1.578181166e-06 pa0 = -2.855530773e-12
+ ags = 4.177671586e-01 lags = -5.195777995e-08 wags = -1.557031386e-06 pags = 5.190163022e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.984076421e-03 lketa = 9.781949960e-09 wketa = 4.996770669e-07 pketa = -9.771378803e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.765408299e-01 lpclm = 2.522435828e-08 wpclm = 1.046784548e-06 ppclm = -2.519709882e-12
+ pdiblc1 = 4.137574096e-01 lpdiblc1 = -4.777106666e-08 wpdiblc1 = -2.373173546e-06 ppdiblc1 = 4.771944142e-12
+ pdiblc2 = 2.902975442e-03 lpdiblc2 = 1.206582560e-10 wpdiblc2 = 1.874078111e-08 ppdiblc2 = -1.205278630e-14
+ pdiblcb = -2.314169863e-02 lpdiblcb = -3.736646369e-09 wpdiblcb = -1.856293136e-07 ppdiblcb = 3.732608250e-13
+ drout = 5.375281665e-01 ldrout = 4.518604815e-08 wdrout = 2.244754862e-06 pdrout = -4.513721650e-12
+ pscbe1 = 7.596311908e+08 lpscbe1 = 8.117303628e+01 wpscbe1 = 4.032518339e+03 ppscbe1 = -8.108531420e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.255049513e-07 lalpha0 = -3.931186189e-13 walpha0 = -1.952936730e-11 palpha0 = 3.926937835e-17
+ alpha1 = 8.525468078e-01 lalpha1 = -5.121085457e-09 walpha1 = -2.544055510e-07 palpha1 = 5.115551203e-13
+ beta0 = 1.406763974e+01 lbeta0 = -4.175190849e-07 wbeta0 = -2.074153492e-05 pbeta0 = 4.170678804e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.106429615e-01 lkt1 = -7.725308033e-09 wkt1 = -4.492178678e-07 pkt1 = 7.716959447e-13
+ kt2 = -4.493098135e-02 lkt2 = -3.021710482e-09 wkt2 = -1.502150554e-07 pkt2 = 3.018444980e-13
+ at = 1.379939085e+05 lat = 7.768084158e-03 wat = 2.003923556e-01 pat = -7.759689345e-7
+ ute = -1.801420659e+00 lute = -1.247256600e-07 wute = -5.172338457e-06 pute = 1.245908715e-11
+ ua1 = 2.851161315e-10 lua1 = -2.588958578e-16 wua1 = -1.059415188e-14 pua1 = 2.586160742e-20
+ ub1 = -4.357671071e-19 lub1 = 1.359264559e-25 wub1 = 5.393875348e-24 pub1 = -1.357795629e-29
+ uc1 = 3.136246856e-11 luc1 = -2.926732120e-18 wuc1 = -1.003963420e-16 puc1 = 2.923569259e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.5 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.171853786e-01 lvth0 = 4.730281984e-09 wvth0 = 6.264239100e-08 pvth0 = 1.740423273e-13
+ k1 = 5.402511595e-01 lk1 = 7.348844679e-09 wk1 = 9.882211729e-07 pk1 = -7.472983274e-13
+ k2 = -2.611597326e-02 lk2 = -5.006548271e-09 wk2 = -4.201058587e-07 pk2 = 3.081479688e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 9.216734667e-01 ldsub = -3.431026432e-07 wdsub = -5.514221115e-06 pdsub = 3.328942642e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.009799929e-01 lvoff = 7.459654747e-10 wvoff = -3.942667057e-08 pvoff = -1.022192820e-13
+ nfactor = 2.651060692e+00 lnfactor = 5.810659875e-08 wnfactor = -1.378147636e-06 pnfactor = 1.012636380e-12
+ eta0 = 2.098785464e-01 leta0 = -1.254765336e-07 weta0 = -4.861098268e-06 peta0 = 4.333868896e-12
+ etab = -1.514243402e-01 letab = 7.708256352e-08 wetab = 1.041452527e-06 petab = -5.312477862e-13
+ u0 = 3.290551512e-02 lu0 = -1.605195596e-09 wu0 = -3.838977123e-08 pu0 = 6.325351285e-16
+ ua = -5.246086823e-10 lua = -1.785475059e-16 wua = -5.159390749e-15 pua = 4.445976670e-23
+ ub = 1.302653397e-18 lub = 1.438810395e-25 wub = 5.412114832e-24 pub = -5.208802570e-31
+ uc = 8.743480464e-12 luc = 3.317321575e-17 wuc = 2.052528342e-16 puc = -7.294601488e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.011565249e+04 lvsat = -1.637493983e-03 wvsat = -1.155275070e-02 pvsat = 1.635724376e-7
+ a0 = 1.285218759e+00 la0 = -7.136336130e-09 wa0 = -4.131210800e-06 pa0 = 2.915442695e-12
+ ags = 2.421556360e-01 lags = 1.255478885e-07 wags = 1.867376187e-06 pags = 1.728819788e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.552025509e-03 lketa = -8.677943660e-10 wketa = -7.420484664e-07 pketa = 2.779809047e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.430483739e-01 lpclm = -4.200053613e-08 wpclm = -2.752738181e-06 ppclm = 1.320794500e-12
+ pdiblc1 = 3.886654915e-01 lpdiblc1 = -2.240850714e-08 wpdiblc1 = 1.333066290e-07 ppdiblc1 = 2.238429072e-12
+ pdiblc2 = 1.088563979e-03 lpdiblc2 = 1.954639961e-09 wpdiblc2 = 2.427070621e-08 ppdiblc2 = -1.764235717e-14
+ pdiblcb = -2.871660273e-02 lpdiblcb = 1.898388643e-09 wpdiblcb = 3.712586273e-07 ppdiblcb = -1.896337092e-13
+ drout = 6.003068905e-01 ldrout = -1.826980710e-08 wdrout = -4.026333161e-06 pdrout = 1.825006329e-12
+ pscbe1 = 8.626304063e+08 lpscbe1 = -2.293712868e+01 wpscbe1 = -6.256272284e+03 ppscbe1 = 2.291234098e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 9.095149961e-08 lalpha0 = -2.571138738e-13 walpha0 = -6.088563054e-12 palpha0 = 2.568360159e-17
+ alpha1 = 8.449063844e-01 lalpha1 = 2.601747532e-09 walpha1 = 5.088111020e-07 palpha1 = -2.598935876e-13
+ beta0 = 1.381870533e+01 lbeta0 = -1.658996662e-07 wbeta0 = 4.125004454e-06 pbeta0 = 1.657203817e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.088932651e-01 lkt1 = -9.493876666e-09 wkt1 = 2.780952962e-07 pkt1 = 3.653798084e-14
+ kt2 = -4.863894634e-02 lkt2 = 7.262486249e-10 wkt2 = 2.215918350e-07 pkt2 = -7.397270157e-14
+ at = 1.724245120e+05 lat = -2.703388781e-02 wat = -6.816543185e-01 pat = 1.155914950e-7
+ ute = -2.117471039e+00 lute = 1.947336395e-07 wute = 1.228547208e-05 pute = -5.187023334e-12
+ ua1 = -3.889710299e-10 lua1 = 4.224620078e-16 wua1 = 2.548682287e-14 pua1 = -1.060853673e-20
+ ub1 = -7.957208323e-20 lub1 = -2.241104874e-25 wub1 = -1.145746394e-23 pub1 = 3.455141541e-30
+ uc1 = 1.652876450e-11 luc1 = 1.206696827e-17 wuc1 = 7.610674947e-16 puc1 = -5.783986598e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.6 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.227670599e-01 lvth0 = 1.879237320e-09 wvth0 = 7.708900208e-07 pvth0 = -1.877206466e-13
+ k1 = 5.759751139e-01 lk1 = -1.089845111e-08 wk1 = -2.606171909e-06 pk1 = 1.088667337e-12
+ k2 = -4.265052859e-02 lk2 = 3.439071106e-09 wk2 = 8.557384789e-07 pk2 = -3.435354570e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.625148754e-01 ldsub = -6.413663034e-09 wdsub = -2.512157659e-07 pdsub = 6.406731917e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.001421779e-01 lvoff = 3.180212539e-10 wvoff = -1.773543439e-07 pvoff = -3.176775747e-14
+ nfactor = 2.789046350e+00 lnfactor = -1.237454362e-08 wnfactor = -1.815670767e-06 pnfactor = 1.236117070e-12
+ eta0 = -3.577527649e-02 weta0 = 3.623607453e-6
+ etab = -5.592675218e-04 letab = 2.279648880e-11 wetab = 5.851314939e-09 petab = -2.277185309e-15
+ u0 = 2.914241571e-02 lu0 = 3.169428958e-10 wu0 = 2.483156476e-08 pu0 = -3.166003820e-14
+ ua = -9.139636730e-10 lua = 2.032957240e-17 wua = -1.096593353e-15 pua = -2.030760264e-21
+ ub = 1.603607069e-18 lub = -9.841882920e-27 wub = 2.467623486e-24 pub = 9.831246994e-31
+ uc = 7.383107134e-11 luc = -7.261444363e-20 wuc = 4.824067653e-17 puc = 7.253597065e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.068210421e+04 lvsat = -1.926829592e-03 wvsat = -6.813670751e-02 pvsat = 1.924747306e-7
+ a0 = 1.271247476e+00 wa0 = 1.576546842e-6
+ ags = 3.928289067e-01 lags = 4.858609127e-08 wags = 1.475374800e-05 pags = -4.853358525e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.481237729e-04 lketa = 4.622421863e-10 wketa = -1.074281562e-07 pketa = -4.617426504e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.511882494e-01 lpclm = 4.920329430e-09 wpclm = 7.953146481e-07 ppclm = -4.915012128e-13
+ pdiblc1 = 2.766248118e-01 lpdiblc1 = 3.482030347e-08 wpdiblc1 = 1.132526659e-05 ppdiblc1 = -3.478267387e-12
+ pdiblc2 = 4.846842543e-03 lpdiblc2 = 3.496388620e-11 wpdiblc2 = -3.431202270e-09 ppdiblc2 = -3.492610142e-15
+ pdiblcb = -4.046081186e-02 lpdiblcb = 7.897166246e-09 wpdiblcb = 1.544410367e-06 ppdiblcb = -7.888631936e-13
+ drout = 6.032873391e-01 ldrout = -1.979217853e-08 wdrout = -4.324055932e-06 pdrout = 1.977078952e-12
+ pscbe1 = 8.362144241e+08 lpscbe1 = -9.444214796e+00 wpscbe1 = -3.617528787e+03 ppscbe1 = 9.434008622e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.721592095e-07 lalpha0 = 1.326723929e-13 walpha0 = 7.014004001e-11 palpha0 = -1.325290165e-17
+ alpha1 = 0.85
+ beta0 = 1.351919086e+01 lbeta0 = -1.291186681e-08 wbeta0 = 3.404408377e-05 pbeta0 = 1.289791322e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.286328252e-01 lkt1 = 5.888142947e-10 wkt1 = 4.647796970e-07 pkt1 = -5.881779749e-14
+ kt2 = -4.751653897e-02 lkt2 = 1.529386538e-10 wkt2 = 1.066799855e-07 pkt2 = -1.527733760e-14
+ at = 1.173723186e+05 lat = 1.086001837e-03 wat = -2.429690048e-01 pat = -1.084828216e-7
+ ute = -1.693075960e+00 lute = -2.204142494e-08 wute = -2.180045486e-06 pute = 2.201760521e-12
+ ua1 = 4.642273863e-10 lua1 = -1.333979846e-17 wua1 = 2.108979768e-15 pua1 = 1.332538240e-21
+ ub1 = -4.849345502e-19 lub1 = -1.705701435e-26 wub1 = -8.028858962e-24 pub1 = 1.703858118e-30
+ uc1 = 4.817616651e-11 luc1 = -4.098081613e-18 wuc1 = -1.172744218e-15 puc1 = 4.093652898e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.7 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.223204654e-01 lvth0 = 1.995702910e-09 wvth0 = 8.155012068e-07 pvth0 = -1.993546193e-13
+ k1 = 5.594265456e-01 lk1 = -6.582816168e-09 wk1 = -9.531034461e-07 pk1 = 6.575702251e-13
+ k2 = -3.909373375e-02 lk2 = 2.511508806e-09 wk2 = 5.004433705e-07 pk2 = -2.508794669e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.058087301e-01 ldsub = 8.374505792e-09 wdsub = 5.413270651e-06 pdsub = -8.365455631e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.014532215e-01 lvoff = 6.599230758e-10 wvoff = -4.639166355e-08 pvoff = -6.592099101e-14
+ nfactor = 2.754218570e+00 lnfactor = -3.291946142e-09 wnfactor = 1.663343481e-06 pnfactor = 3.288388602e-13
+ eta0 = -1.284871776e-01 leta0 = 2.417796585e-08 weta0 = 1.288477838e-05 peta0 = -2.415183720e-12
+ etab = -6.019751828e-03 letab = 1.446814349e-09 wetab = 5.513096419e-07 petab = -1.445250806e-13
+ u0 = 3.359495311e-02 lu0 = -8.442165210e-10 wu0 = -4.199409978e-07 pu0 = 8.433041931e-14
+ ua = -5.614905365e-10 lua = -7.159048698e-17 wua = -3.630581594e-14 pua = 7.151312057e-21
+ ub = 1.389162684e-18 lub = 4.608221042e-26 wub = 2.388888739e-23 pub = -4.603241030e-30
+ uc = 7.391841099e-11 luc = -9.539139970e-20 wuc = 3.951615088e-17 puc = 9.528831212e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.363106444e+04 lvsat = -8.801713357e-05 wvsat = 6.362052782e-01 pvsat = 8.792201522e-9
+ a0 = 1.271247476e+00 wa0 = 1.576546842e-6
+ ags = 8.276643286e-01 lags = -6.481289906e-08 wags = -2.868280239e-05 pags = 6.474285706e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.581967936e-03 lketa = 3.615850247e-11 wketa = -2.706360062e-07 pketa = -3.611942670e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.446950564e-01 lpclm = 6.613663250e-09 wpclm = 1.443932238e-06 ppclm = -6.606515997e-13
+ pdiblc1 = 4.619969338e-01 lpdiblc1 = -1.352215071e-08 wpdiblc1 = -7.191912812e-06 ppdiblc1 = 1.350753760e-12
+ pdiblc2 = 6.251297878e-03 lpdiblc2 = -3.312984028e-10 wpdiblc2 = -1.437249591e-07 ppdiblc2 = 3.309403752e-14
+ pdiblcb = 1.782452985e-02 lpdiblcb = -7.302834878e-09 wpdiblcb = -4.277825024e-06 ppdiblcb = 7.294942850e-13
+ drout = 4.702130150e-01 ldrout = 1.491174215e-08 wdrout = 8.968995400e-06 pdrout = -1.489562733e-12
+ pscbe1 = 7.991711766e+08 lpscbe1 = 2.161455343e-01 wpscbe1 = 8.279276883e+01 ppscbe1 = -2.159119501e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.946638415e-07 lalpha0 = 1.385412859e-13 walpha0 = 7.238807117e-11 palpha0 = -1.383915671e-17
+ alpha1 = 9.188950814e-01 lalpha1 = -1.796687269e-08 walpha1 = -6.882062782e-06 palpha1 = 1.794745625e-12
+ beta0 = 1.263611164e+01 lbeta0 = 2.173828308e-07 wbeta0 = 1.222565732e-04 pbeta0 = -2.171479095e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.198038924e-01 lkt1 = -1.713647765e-09 wkt1 = -4.171594542e-07 pkt1 = 1.711795860e-13
+ kt2 = -4.616455406e-02 lkt2 = -1.996400831e-10 wkt2 = -2.837239922e-08 pkt2 = 1.994243361e-14
+ at = 1.235649369e+05 lat = -5.289463121e-04 wat = -8.615616081e-01 pat = 5.283746904e-8
+ ute = -1.970598865e+00 lute = 5.033266315e-08 wute = 2.554225359e-05 pute = -5.027826965e-12
+ ua1 = 5.995254285e-12 lua1 = 1.061607263e-16 wua1 = 4.788267274e-14 pua1 = -1.060460006e-20
+ ub1 = -2.101392518e-19 lub1 = -8.871978104e-26 wub1 = -3.547869222e-23 pub1 = 8.862390335e-30
+ uc1 = 4.085764812e-11 luc1 = -2.189514478e-18 wuc1 = -4.416832776e-16 puc1 = 2.187148314e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.8 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.268831981e-01 lvth0 = 1.125197404e-09 wvth0 = 3.597210303e-07 pvth0 = -1.123981426e-13
+ k1 = 5.312785764e-01 lk1 = -1.212577708e-09 wk1 = 1.858651584e-06 pk1 = 1.211267300e-13
+ k2 = -3.087042946e-02 lk2 = 9.426174735e-10 wk2 = -3.209983826e-07 pk2 = -9.415988056e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.209432474e-01 ldsub = 5.487051776e-09 wdsub = 3.901454479e-06 pdsub = -5.481122029e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 3.255239980e-03 lcdscd = 4.091902473e-10 wcdscd = 2.142442546e-07 pcdscd = -4.087480436e-14
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.230164554e-01 lvoff = 4.773886218e-09 wvoff = 2.107601431e-06 pvoff = -4.768727175e-13
+ nfactor = 1.877145382e+00 lnfactor = 1.640413391e-07 wnfactor = 8.927587873e-05 pnfactor = -1.638640629e-11
+ eta0 = -1.375413602e-02 leta0 = 2.288507773e-09 weta0 = 1.423873186e-06 peta0 = -2.286034628e-13
+ etab = -4.088343487e-03 letab = 1.078328677e-09 wetab = 3.583775313e-07 petab = -1.077163349e-13
+ u0 = 2.412533861e-02 lu0 = 9.624533496e-10 wu0 = 5.259970892e-07 pu0 = -9.614132455e-14
+ ua = -1.561762283e-09 lua = 1.192473585e-16 wua = 6.361326137e-14 pua = -1.191184903e-20
+ ub = 2.182599896e-18 lub = -1.052945015e-25 wub = -5.536908863e-23 pub = 1.051807118e-29
+ uc = 6.020391540e-11 luc = 2.521142355e-18 wuc = 1.409483611e-15 puc = -2.518417807e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.953013081e+04 lvsat = -1.213476411e-03 wvsat = 4.693614096e-02 pvsat = 1.212165031e-7
+ a0 = 1.271247476e+00 wa0 = 1.576546842e-6
+ ags = 4.879491552e-01 wags = 5.252002603e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.729722354e-02 lketa = -4.679166254e-09 wketa = -2.739490639e-06 pketa = 4.674109572e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.329144285e-01 lpclm = 8.861242133e-09 wpclm = 2.620721924e-06 ppclm = -8.851665966e-13
+ pdiblc1 = 3.958216889e-01 lpdiblc1 = -8.968404512e-10 wpdiblc1 = -5.815397536e-07 ppdiblc1 = 8.958712537e-14
+ pdiblc2 = 4.801725630e-03 lpdiblc2 = -5.474031191e-11 wpdiblc2 = 1.075613326e-09 ppdiblc2 = 5.468115515e-15
+ pdiblcb = 1.384183335e-02 lpdiblcb = -6.542992142e-09 wpdiblcb = -3.879985776e-06 ppdiblcb = 6.535921262e-13
+ drout = 4.767543002e-01 ldrout = 1.366375651e-08 wdrout = 8.315573786e-06 pdrout = -1.364899037e-12
+ pscbe1 = 7.981748633e+08 lpscbe1 = 4.062281646e-01 wpscbe1 = 1.823164298e+02 ppscbe1 = -4.057891619e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.951900711e-08 lalpha0 = -1.530523077e-15 walpha0 = -9.508720107e-13 palpha0 = 1.528869071e-19
+ alpha1 = 6.892448102e-01 lalpha1 = 2.584718395e-08 walpha1 = 1.605814649e-05 palpha1 = -2.581925142e-12
+ beta0 = 1.332273551e+01 lbeta0 = 8.638460776e-08 wbeta0 = 5.366838757e-05 pbeta0 = -8.629125364e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.114258703e-01 lkt1 = -3.312057091e-09 wkt1 = -1.254056269e-06 pkt1 = 3.308477817e-13
+ kt2 = -4.453891522e-02 lkt2 = -5.097892149e-10 wkt2 = -1.907606037e-07 pkt2 = 5.092382959e-14
+ at = 1.195066423e+05 lat = 2.453194799e-04 wat = -4.561707207e-01 pat = -2.450543680e-8
+ ute = -9.821497330e-01 lute = -1.382495928e-07 wute = -7.319583984e-05 pute = 1.381001893e-11
+ ua1 = 1.571650889e-09 lua1 = -1.925444496e-16 wua1 = -1.085136935e-13 pua1 = 1.923363707e-20
+ ub1 = -1.253525650e-18 lub1 = 1.103437364e-25 wub1 = 6.874719095e-23 pub1 = -1.102244901e-29
+ uc1 = 4.017607318e-11 luc1 = -2.059479521e-18 wuc1 = -3.735994396e-16 puc1 = 2.057253882e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.9 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.188593681e-01 lvth0 = -2.772767157e-07 wvth0 = -1.910766174e-08 pvth0 = 1.910972270e-12
+ k1 = 5.418064353e-01 lk1 = -9.408868149e-08 wk1 = -6.483828602e-09 pk1 = 6.484527948e-13
+ k2 = -2.769247282e-02 lk2 = 9.842879788e-08 wk2 = 6.782914213e-09 pk2 = -6.783645819e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.045417318e-01 lvoff = -7.269465504e-08 wvoff = -5.009525865e-09 pvoff = 5.010066193e-13
+ nfactor = 2.550155693e+00 lnfactor = 1.343888008e-05 wnfactor = 9.260985874e-07 pnfactor = -9.261984764e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.149477126e-02 lu0 = -3.267478013e-09 wu0 = -2.251680762e-10 pu0 = 2.251923628e-14
+ ua = -7.366463064e-10 lua = -2.131506240e-15 wua = -1.468861175e-16 pua = 1.469019606e-20
+ ub = 1.537372114e-18 lub = 3.312145784e-24 wub = 2.282462165e-25 pub = -2.282708352e-29
+ uc = 4.773753148e-11 luc = 1.504630793e-16 wuc = 1.036869474e-17 puc = -1.036981311e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.376452071e+00 la0 = -7.001826012e-07 wa0 = -4.825090441e-08 pa0 = 4.825610875e-12
+ ags = 3.811550339e-01 lags = -1.130155785e-07 wags = -7.788116792e-09 pags = 7.788956818e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 8.180254810e-25 lb1 = 1.289455985e-28 wb1 = 8.885884532e-30 pb1 = -8.886842964e-34
+ keta = -7.199184736e-03 lketa = -1.595587346e-07 wketa = -1.099549351e-08 pketa = 1.099667949e-12
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.725335471e-02 lpclm = -3.094069161e-06 wpclm = -2.132181449e-07 ppclm = 2.132411426e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.147018095e-03 lpdiblc2 = -7.356732866e-09 wpdiblc2 = -5.069663451e-10 ppdiblc2 = 5.070210265e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.178768667e+08 lpscbe1 = 3.680126221e+03 wpscbe1 = 2.536044429e+02 ppscbe1 = -2.536317966e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.199864079e-01 lkt1 = 6.957158242e-07 wkt1 = 4.794309037e-08 pkt1 = -4.794826152e-12
+ kt2 = -4.543335553e-02 lkt2 = 1.200314779e-08 wkt2 = 8.271595661e-10 pkt2 = -8.272487835e-14
+ at = 140000.0
+ ute = -1.856411036e+00 lute = 4.301567497e-06 wute = 2.964291340e-07 pute = -2.964611068e-11
+ ua1 = 3.044858563e-10 lua1 = 7.154185942e-15 wua1 = 4.930084544e-16 pua1 = -4.930616303e-20
+ ub1 = -5.528820975e-19 lub1 = -8.674725804e-24 wub1 = -5.977917258e-25 pub1 = 5.978562036e-29
+ uc1 = 1.656219400e-11 luc1 = -7.325600042e-17 wuc1 = -5.048209235e-18 puc1 = 5.048753735e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.10 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.050030051e-01 wvth0 = 7.638945015e-8
+ k1 = 5.371045370e-01 wk1 = 2.592133503e-8
+ k2 = -2.277368563e-02 wk2 = -2.711703264e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.081745054e-01 wvoff = 2.002730274e-8
+ nfactor = 3.221737513e+00 wnfactor = -3.702397647e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.133148542e-02 wu0 = 9.001868339e-10
+ ua = -8.431641733e-10 wua = 5.872277781e-16
+ ub = 1.702890140e-18 wub = -9.124927588e-25
+ uc = 5.525663039e-11 wuc = -4.145242368e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.341461811e+00 wa0 = 1.928995869e-7
+ ags = 3.755073008e-01 wags = 3.113567570e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 7.261830261e-24 wb1 = -3.552437983e-29
+ keta = -1.517282128e-02 wketa = 4.395826736e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.736671676e-02 wpclm = 8.524128735e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.779379719e-03 wpdiblc2 = 2.026772342e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.017839967e+08 wpscbe1 = -1.013870991e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.852193666e-01 wkt1 = -1.916689944e-7
+ kt2 = -4.483352163e-02 wkt2 = -3.306854877e-9
+ at = 140000.0
+ ute = -1.641448590e+00 wute = -1.185077424e-6
+ ua1 = 6.620023447e-10 wua1 = -1.970970873e-15
+ ub1 = -9.863845998e-19 wub1 = 2.389878042e-24
+ uc1 = 1.290136826e-11 wuc1 = 2.018195281e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.11 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.865892412e-01 lvth0 = 1.475087222e-07 wvth0 = 1.471195825e-07 pvth0 = -5.666039541e-13
+ k1 = 5.246957231e-01 lk1 = 9.940435247e-08 wk1 = 4.822739943e-08 pk1 = -1.786891084e-13
+ k2 = -1.122526934e-02 lk2 = -9.251189154e-08 wk2 = -6.859979467e-08 pk2 = 3.323095293e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.176113977e-01 lvoff = 7.559692437e-08 wvoff = 6.005283304e-08 pvoff = -3.206359578e-13
+ nfactor = 3.787202708e+00 lnfactor = -4.529820674e-06 wnfactor = -7.739483276e-06 pnfactor = 3.234022904e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.189532637e-02 lu0 = -4.516809250e-09 wu0 = 6.263600579e-10 pu0 = 2.193567704e-15
+ ua = -8.804820293e-10 lua = 2.989453581e-16 wua = 8.064207034e-16 pua = -1.755907617e-21
+ ub = 1.877153765e-18 lub = -1.395988610e-24 wub = -1.585058649e-24 pub = 5.387781416e-30
+ uc = 1.749290886e-10 luc = -9.586704525e-16 wuc = -8.223658220e-16 puc = 6.255730119e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.769452386e+00 la0 = -3.428540902e-06 wa0 = -2.039645614e-06 pa0 = 1.788444184e-11
+ ags = 4.476107193e-01 lags = -5.776050552e-07 wags = -6.188986654e-07 pags = 5.207285999e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.454324205e-23 lb1 = -5.832983160e-29 wb1 = -7.114455115e-29 pb1 = 2.853455697e-34
+ keta = -2.844591055e-02 lketa = 1.063278777e-07 wketa = 8.835622306e-08 pketa = -3.556625219e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.020884212e+00 lpclm = 7.398101022e-06 wpclm = 3.342478635e-06 ppclm = -1.994738394e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.818096188e-03 lpdiblc2 = -3.101493542e-10 wpdiblc2 = 1.641582583e-09 ppdiblc2 = 3.085672732e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.001221352e+09 lpscbe1 = -7.965713764e+02 wpscbe1 = -2.012411431e+03 ppscbe1 = 7.999093778e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.601231753e-01 lkt1 = -2.010402180e-07 wkt1 = -3.500490494e-07 pkt1 = 1.268748728e-12
+ kt2 = -3.219755090e-02 lkt2 = -1.012240574e-07 wkt2 = -8.264351494e-08 pkt2 = 6.355490057e-13
+ at = 140000.0
+ ute = -1.123537024e+00 lute = -4.148878724e-06 wute = -4.479450180e-06 pute = 2.639051515e-11
+ ua1 = 1.912795055e-09 lua1 = -1.001983273e-14 wua1 = -9.230253929e-15 pua1 = 5.815256307e-20
+ ub1 = -2.186713527e-18 lub1 = 9.615578161e-24 wub1 = 8.880586807e-24 pub1 = -5.199567891e-29
+ uc1 = -2.771450635e-11 luc1 = 3.253650797e-16 wuc1 = 1.997098526e-16 puc1 = -1.438159586e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.12 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.238910272e-01 lvth0 = -2.100759086e-09 wvth0 = -4.119398830e-08 pvth0 = 1.886814793e-13
+ k1 = 5.756552523e-01 lk1 = -1.049834137e-07 wk1 = -1.758356650e-07 pk1 = 7.199798934e-13
+ k2 = -4.225743877e-02 lk2 = 3.195149914e-08 wk2 = 8.205363029e-08 pk2 = -2.719291184e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -8.871247706e-02 lvoff = -4.031046194e-08 wvoff = -8.729703218e-08 pvoff = 2.703528187e-13
+ nfactor = 2.520055606e+00 lnfactor = 5.524351856e-07 wnfactor = 8.151637335e-07 pnfactor = -1.970629421e-12
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398724195e-01 letab = 2.802433220e-07 wetab = -1.171062741e-11 petab = 4.696882045e-17
+ u0 = 3.207753642e-02 lu0 = -5.247614758e-09 wu0 = 2.885059913e-09 pu0 = -6.865594051e-15
+ ua = -4.011086334e-10 lua = -1.623718747e-15 wua = -1.226352763e-15 pua = 6.397111744e-21
+ ub = 9.744011767e-19 lub = 2.224758832e-24 wub = 2.650668732e-24 pub = -1.160081466e-29
+ uc = -2.093422232e-10 luc = 5.825595450e-16 wuc = 1.520696392e-15 puc = -3.141791005e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 4.153275676e-01 la0 = 2.002563960e-06 wa0 = 5.712583713e-06 pa0 = -1.320809101e-11
+ ags = 1.144642986e-01 lags = 7.585739446e-07 wags = 1.024303754e-06 pags = -1.383247261e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.180386289e-05 lketa = -7.635023608e-09 wketa = -2.629050060e-08 pketa = 1.041609523e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.320634398e-01 lpclm = -3.367547891e-08 wpclm = -1.495708702e-06 ppclm = -5.424499062e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.305949366e-03 lpdiblc2 = 5.754747951e-09 wpdiblc2 = 3.683254340e-10 ppdiblc2 = 8.192434679e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.052422032e+08 lpscbe1 = -1.054094871e+01 wpscbe1 = -3.612890767e+01 ppscbe1 = 7.264750173e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.046064812e-01 lkt1 = -2.262719718e-08 wkt1 = -1.134304931e-08 pkt1 = -8.972855592e-14
+ kt2 = -5.800521569e-02 lkt2 = 2.284963183e-09 wkt2 = 7.983863007e-08 pkt2 = -1.613210674e-14
+ at = 1.682199118e+05 lat = -1.131840272e-01 wat = -2.084646247e-02 pat = 8.361069983e-8
+ ute = -2.533092297e+00 lute = 1.504545829e-06 wute = 3.727476919e-06 pute = -6.525713158e-12
+ ua1 = -1.720323789e-09 lua1 = 4.551829464e-15 wua1 = 1.096817911e-14 pua1 = -2.285902938e-20
+ ub1 = 1.238884608e-18 lub1 = -4.123762879e-24 wub1 = -9.897674307e-24 pub1 = 2.331990787e-29
+ uc1 = 6.694697625e-11 luc1 = -5.430186945e-17 wuc1 = -2.942920936e-16 puc1 = 5.431765036e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.13 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.943497501e-01 lvth0 = 5.730042734e-08 wvth0 = 7.171955536e-08 pvth0 = -3.836349352e-14
+ k1 = 4.320314661e-01 lk1 = 1.838132848e-07 wk1 = 5.771236946e-07 pk1 = -7.940602453e-13
+ k2 = 1.043823076e-02 lk2 = -7.400821541e-08 wk2 = -2.113560778e-07 pk2 = 3.180550150e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.152362433e+00 ldsub = -1.794349887e-06 wdsub = -6.150101207e-06 pdsub = 1.236653740e-11
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.036330347e-01 lvoff = -1.030841350e-08 wvoff = 1.422205481e-07 pvoff = -1.911579184e-13
+ nfactor = 2.908375480e+00 lnfactor = -2.283929821e-07 wnfactor = -1.331454003e-07 pnfactor = -6.378269137e-14
+ eta0 = -6.590106194e-03 leta0 = 1.425668627e-08 weta0 = 3.471429712e-08 peta0 = -6.980302264e-14
+ etab = -9.758147600e-04 letab = 9.519737058e-10 wetab = 1.963530663e-09 petab = -3.924818713e-15
+ u0 = 3.309312078e-02 lu0 = -7.289737565e-09 wu0 = -7.636131088e-10 pu0 = 4.711065784e-16
+ ua = -9.099793181e-10 lua = -6.004886983e-16 wua = 3.509173667e-15 pua = -3.125018505e-21
+ ub = 1.950124731e-18 lub = 2.627875688e-25 wub = -5.890541933e-24 pub = 5.573732167e-30
+ uc = 7.457786857e-11 luc = 1.165699933e-17 wuc = 9.181504903e-17 puc = -2.686164054e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.885541875e+04 lvsat = 1.229486679e-01 wvsat = 2.799890480e-01 pvsat = -5.629980579e-7
+ a0 = 2.455556164e+00 la0 = -2.099899139e-06 wa0 = -6.731274788e-06 pa0 = 1.181384545e-11
+ ags = 9.420035339e-01 lags = -9.054303641e-07 wags = -5.170032837e-06 pags = 1.107223804e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.356607466e-02 lketa = -1.154088874e-07 wketa = 8.236954313e-08 pketa = -1.143311424e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.101756931e+00 lpclm = -5.759713759e-07 wpclm = -2.572969108e-06 ppclm = 1.623690236e-12
+ pdiblc1 = -2.053601678e-01 lpdiblc1 = 1.197141890e-06 wpdiblc1 = 1.893742697e-06 ppdiblc1 = -3.807911303e-12
+ pdiblc2 = 6.892558304e-03 lpdiblc2 = -5.478727089e-09 wpdiblc2 = -8.755152680e-09 ppdiblc2 = 2.653779674e-14
+ pdiblcb = -4.984180035e-02 lpdiblcb = 4.995154436e-08 wpdiblcb = -1.614028203e-09 ppdiblcb = 3.245465313e-15
+ drout = 8.632358000e-01 ldrout = -6.097423013e-7
+ pscbe1 = 2.367661598e+09 lpscbe1 = -3.152231995e+03 wpscbe1 = -7.049917884e+03 ppscbe1 = 1.417587618e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.586663671e-07 lalpha0 = -6.608777297e-13 walpha0 = -2.044710672e-11 palpha0 = 4.111475594e-17
+ alpha1 = 8.156332760e-01 lalpha1 = 6.910412749e-8
+ beta0 = 1.174294166e+01 lbeta0 = 4.256951278e-06 wbeta0 = -4.719873801e-06 pbeta0 = 9.490656162e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.617030336e-01 lkt1 = 9.218175103e-08 wkt1 = -9.731532246e-08 pkt1 = 8.314328732e-14
+ kt2 = -8.777548880e-02 lkt2 = 6.214661158e-08 wkt2 = 1.450663766e-07 pkt2 = -1.472911463e-13
+ at = 1.579085934e+05 lat = -9.245017255e-02 wat = 6.314170135e-02 pat = -8.527152414e-8
+ ute = -2.589035663e+00 lute = 1.617035967e-06 wute = 2.558505937e-07 pute = 4.549844548e-13
+ ua1 = -9.103542364e-10 lua1 = 2.923154027e-15 wua1 = -2.355051396e-15 pua1 = 3.931135995e-21
+ ub1 = -3.210116898e-19 lub1 = -9.871452416e-25 wub1 = 4.602988815e-24 pub1 = -5.837822523e-30
+ uc1 = 1.085175074e-11 luc1 = 5.849362467e-17 wuc1 = 4.096213043e-17 puc1 = -1.309479965e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.14 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.324359490e-01 lvth0 = 1.880343073e-08 wvth0 = -4.246350278e-08 pvth0 = 7.705114309e-14
+ k1 = 7.243968413e-01 lk1 = -1.117055434e-07 wk1 = -2.808983443e-07 pk1 = 7.321641923e-14
+ k2 = -1.117546243e-01 lk2 = 4.950261180e-08 wk2 = 1.701099009e-07 pk2 = -6.752545577e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.760407772e+00 ldsub = 1.149837457e-06 wdsub = 1.297050040e-05 pdsub = -6.960299009e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.065630528e-01 lvoff = -7.346792241e-09 wvoff = -9.486017314e-10 pvoff = -4.644454612e-14
+ nfactor = 2.268773401e+00 lnfactor = 4.181078448e-07 wnfactor = 1.256550378e-06 pnfactor = -1.468467728e-12
+ eta0 = -4.853792816e-01 leta0 = 4.982100817e-07 weta0 = -6.942859423e-08 peta0 = 3.546315393e-14
+ etab = 2.505088655e-04 letab = -2.875770464e-10 wetab = -3.880218816e-09 petab = 1.981961448e-15
+ u0 = 2.852315666e-02 lu0 = -2.670481817e-09 wu0 = -8.186854767e-09 pu0 = 7.974415321e-15
+ ua = -1.260373075e-09 lua = -2.463155942e-16 wua = -8.855258609e-17 pua = 5.115128236e-22
+ ub = 2.114752812e-18 lub = 9.638380952e-26 wub = -1.848191152e-25 pub = -1.935325775e-31
+ uc = 8.651100948e-11 luc = -4.048524357e-19 wuc = -3.307156876e-16 puc = 1.584717478e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.818236357e+05 lvsat = -4.177732423e-02 wvsat = -7.125172551e-01 pvsat = 4.402134182e-7
+ a0 = -7.680726914e-01 la0 = 1.158499778e-06 wa0 = 1.001993426e-05 pa0 = -5.118042139e-12
+ ags = -1.183497760e+00 lags = 1.242996587e-06 wags = 1.169288245e-05 pags = -5.972560655e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.287715622e-02 lketa = 2.250602020e-08 wketa = -1.463844231e-07 pketa = 1.168901641e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.454808005e-01 lpclm = 2.895405492e-07 wpclm = -1.272950021e-08 ppclm = -9.641641155e-13
+ pdiblc1 = 6.539326663e-01 lpdiblc1 = 3.285807237e-07 wpdiblc1 = -1.694896701e-06 ppdiblc1 = -1.805648400e-13
+ pdiblc2 = -1.581019058e-03 lpdiblc2 = 3.086246279e-09 wpdiblc2 = 4.266929097e-08 ppdiblc2 = -2.544131096e-14
+ pdiblcb = 2.468360070e-02 lpdiblcb = -2.537768767e-08 wpdiblcb = 3.228056405e-09 ppdiblcb = -1.648846019e-15
+ drout = 1.061865782e+00 ldrout = -8.105147058e-07 wdrout = -7.207365652e-06 pdrout = 7.285104298e-12
+ pscbe1 = -1.493337837e+09 lpscbe1 = 7.504121807e+02 wpscbe1 = 9.980900644e+03 ppscbe1 = -3.038636754e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.164353793e-05 lalpha0 = 2.157864235e-11 walpha0 = 1.437040602e-10 palpha0 = -1.248069455e-16
+ alpha1 = 9.187334480e-01 lalpha1 = -3.510808297e-8
+ beta0 = 7.038229371e-01 lbeta0 = 1.541513793e-05 wbeta0 = 9.451188209e-05 pbeta0 = -9.081141345e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.685231124e-01 lkt1 = -2.003208800e-09 wkt1 = -1.330503908e-10 pkt1 = -1.508719273e-14
+ kt2 = -1.693659162e-02 lkt2 = -9.456353950e-09 wkt2 = 3.101362028e-09 pkt2 = -3.794897042e-15
+ at = 8.077706654e+04 lat = -1.448670502e-02 wat = -5.002635658e-02 pat = 2.911716446e-8
+ ute = -6.535547181e-01 lute = -3.393210752e-07 wute = 2.196260345e-06 pute = -1.506354556e-12
+ ua1 = 2.635044555e-09 lua1 = -6.604854357e-16 wua1 = 4.645513098e-15 pua1 = -3.144936588e-21
+ ub1 = -1.241995230e-18 lub1 = -5.622797294e-26 wub1 = -3.446122658e-24 pub1 = 2.298106667e-30
+ uc1 = 1.553485586e-10 luc1 = -8.756172578e-17 wuc1 = -1.956690866e-16 puc1 = 1.082355248e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.15 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.200995669e-01 lvth0 = -2.597391799e-08 wvth0 = 1.000810017e-07 pvth0 = 4.241405832e-15
+ k1 = 2.473628332e-01 lk1 = 1.319567495e-07 wk1 = -3.413984157e-07 pk1 = 1.041190087e-13
+ k2 = 6.991576078e-02 lk2 = -4.329207752e-08 wk2 = 7.993926712e-08 pk2 = -2.146755842e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.694105324e-01 ldsub = 6.195608480e-08 wdsub = -9.879333645e-07 pdsub = 1.694735387e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.007302728e-01 lvoff = -1.032609460e-08 wvoff = -1.733012334e-07 pvoff = 4.159076517e-14
+ nfactor = 2.938532925e+00 lnfactor = 7.600405702e-08 wnfactor = -2.845922071e-06 pnfactor = 6.270177640e-13
+ eta0 = 0.49
+ etab = -2.414997841e-04 letab = -3.626591627e-11 wetab = 3.661281299e-09 petab = -1.870131230e-15
+ u0 = 2.953985264e-02 lu0 = -3.189795891e-09 wu0 = 2.209245645e-08 pu0 = -7.491832939e-15
+ ua = -1.304151342e-09 lua = -2.239542685e-16 wua = 1.592553528e-15 pua = -3.471726437e-22
+ ub = 1.901068449e-18 lub = 2.055307907e-25 wub = 4.175398844e-25 pub = -5.012091215e-31
+ uc = -7.331682434e-12 luc = 4.752868080e-17 wuc = 6.076088565e-16 puc = -3.208112929e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.168760594e+04 lvsat = 4.512577789e-02 wvsat = 4.073686830e-01 pvsat = -1.318086406e-7
+ a0 = 1.5
+ ags = 2.533556992e+00 lags = -6.556229419e-07 wags = -4.396182092e-12 pags = 2.245508265e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.321862732e-02 lketa = -7.966721141e-09 wketa = 5.912744897e-08 pketa = 1.191757704e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.264088925e+00 lpclm = -2.307502202e-07 wpclm = -4.117948330e-06 ppclm = 1.132724189e-12
+ pdiblc1 = 3.500271335e+00 lpdiblc1 = -1.125289220e-06 wpdiblc1 = -1.089188604e-05 ppdiblc1 = 4.517128559e-12
+ pdiblc2 = 6.445527389e-03 lpdiblc2 = -1.013601275e-09 wpdiblc2 = -1.444922952e-08 ppdiblc2 = 3.734029647e-15
+ pdiblcb = 6.939277514e-01 lpdiblcb = -3.672182304e-07 wpdiblcb = -3.516945673e-06 ppdiblcb = 1.796406612e-12
+ drout = -2.115658123e+00 ldrout = 8.125200193e-07 wdrout = 1.441473130e-05 pdrout = -3.759160118e-12
+ pscbe1 = -8.839707193e+08 lpscbe1 = 4.391559880e+02 wpscbe1 = 8.237870249e+03 ppscbe1 = -2.148321231e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.408558481e-05 lalpha0 = -1.199487334e-11 walpha0 = -2.383272882e-10 palpha0 = 7.032931888e-17
+ alpha1 = 0.85
+ beta0 = 4.385311210e+01 lbeta0 = -6.624914882e-06 wbeta0 = -1.750152387e-04 pbeta0 = 4.685926649e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.062179859e-01 lkt1 = -3.382779518e-08 wkt1 = -3.788950514e-07 pkt1 = 1.783791347e-13
+ kt2 = 3.728318971e-03 lkt2 = -2.001170097e-08 wkt2 = -2.464960908e-07 pkt2 = 1.236959875e-13
+ at = 8.326673287e+04 lat = -1.575839172e-02 wat = -7.915627080e-03 pat = 7.607593381e-9
+ ute = -1.207134136e+00 lute = -5.656045848e-08 wute = -5.529123494e-06 pute = 2.439663353e-12
+ ua1 = 1.794695167e-09 lua1 = -2.312467333e-16 wua1 = -7.060513702e-15 pua1 = 2.834338018e-21
+ ub1 = -2.211127900e-18 lub1 = 4.387914272e-25 wub1 = 3.867948226e-24 pub1 = -1.437818344e-30
+ uc1 = -1.537784305e-10 luc1 = 7.033601246e-17 wuc1 = 2.191131311e-16 puc1 = -1.036294250e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.16 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.773691330e-01 lvth0 = -1.483041907e-08 wvth0 = 4.361095333e-07 pvth0 = -8.339013080e-14
+ k1 = 3.929471458e-01 lk1 = 9.399039896e-08 wk1 = 1.942612567e-07 pk1 = -3.557353461e-14
+ k2 = 5.258147608e-02 lk2 = -3.877153875e-08 wk2 = -1.313759417e-07 pk2 = 3.364048963e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.149386476e+00 ldsub = -1.414507217e-07 wdsub = -1.089803013e-06 pdsub = 1.960397170e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -4.391585505e-02 lvoff = -2.514249935e-08 wvoff = -4.429352804e-07 pvoff = 1.119075498e-13
+ nfactor = 4.317577045e+00 lnfactor = -2.836313430e-07 wnfactor = -9.111216819e-06 pnfactor = 2.260918920e-12
+ eta0 = 1.785091854e+00 leta0 = -3.377418242e-07 weta0 = -3.034781852e-07 peta0 = 7.914286201e-14
+ etab = 9.694732365e-02 letab = -2.538175042e-08 wetab = -1.583324405e-07 petab = 4.037556351e-14
+ u0 = -3.158093251e-02 lu0 = 1.274964919e-08 wu0 = 2.924677390e-08 pu0 = -9.357578770e-15
+ ua = -5.801454442e-09 lua = 9.488794177e-16 wua = -1.923410210e-16 pua = 1.183028660e-22
+ ub = 4.365278260e-18 lub = -4.371006291e-25 wub = 3.377701223e-24 pub = -1.273177756e-30
+ uc = 3.824859231e-10 luc = -5.413029328e-17 wuc = -2.087110160e-15 puc = 3.819337006e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.305653097e+05 lvsat = 1.412413704e-02 wvsat = 2.438183315e-01 pvsat = -8.915699862e-8
+ a0 = 1.5
+ ags = -3.334132116e+00 lags = 8.745882298e-07 wags = 1.570065032e-11 pags = -2.995464273e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.252174902e-01 lketa = 1.863315431e-08 wketa = 6.101491687e-07 pketa = -1.317811732e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.344731062e+00 lpclm = -2.517805605e-07 wpclm = -4.069861508e-06 ppclm = 1.120183820e-12
+ pdiblc1 = -4.053430367e+00 lpdiblc1 = 8.446104324e-07 wpdiblc1 = 2.392810509e-05 ppdiblc1 = -4.563437650e-12
+ pdiblc2 = -1.144466001e-02 lpdiblc2 = 3.651909135e-09 wpdiblc2 = -2.176562067e-08 ppdiblc2 = 5.642042029e-15
+ pdiblcb = -2.557604613e+00 lpdiblcb = 4.807358888e-07 wpdiblcb = 1.347185750e-05 ppdiblcb = -2.634035412e-12
+ drout = 2.345302393e+00 ldrout = -3.508360297e-07 wdrout = -3.953993084e-06 pdrout = 1.031146040e-12
+ pscbe1 = 8.224207200e+08 lpscbe1 = -5.847009874e+00 wpscbe1 = -7.744150286e+01 ppscbe1 = 2.019565977e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.292487415e-06 lalpha0 = -1.617390645e-12 walpha0 = 3.801696384e-11 palpha0 = -1.737393242e-18
+ alpha1 = -3.544460907e+00 lalpha1 = 1.146013882e-06 walpha1 = 2.387908318e-05 palpha1 = -6.227330586e-12
+ beta0 = 5.046385996e+01 lbeta0 = -8.348905373e-06 wbeta0 = -1.384496959e-04 pbeta0 = 3.732348484e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.365837245e-01 lkt1 = 7.840556432e-08 wkt1 = 1.766065607e-06 pkt1 = -3.809965756e-13
+ kt2 = -1.719377854e-01 lkt2 = 2.579955974e-08 wkt2 = 8.384481588e-07 pkt2 = -1.592422836e-13
+ at = 4.137853949e+04 lat = -4.834537323e-03 wat = -2.951385460e-01 pat = 8.251130951e-8
+ ute = -3.947397095e-01 lute = -2.684215515e-07 wute = 1.468153945e-05 pute = -2.830994593e-12
+ ua1 = 4.987087401e-09 lua1 = -1.063777934e-15 wua1 = 1.355332439e-14 pua1 = -2.541462362e-21
+ ub1 = -5.369234270e-18 lub1 = 1.262381355e-24 wub1 = 7.743982681e-26 pub1 = -4.493068204e-31
+ uc1 = -1.445876184e-10 luc1 = 6.793917735e-17 wuc1 = 8.363928891e-16 puc1 = -2.646073440e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.17 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.090196161e-01 lvth0 = -1.790288133e-09 wvth0 = 4.828356227e-07 pvth0 = -9.230481450e-14
+ k1 = 7.799027841e-01 lk1 = 2.016468055e-08 wk1 = 1.451504503e-07 pk1 = -2.620388030e-14
+ k2 = 2.244796591e-03 lk2 = -2.916800502e-08 wk2 = -5.492262687e-07 pk2 = 1.133604821e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.710797545e+00 ldsub = -2.485600938e-07 wdsub = -6.366520028e-06 pdsub = 1.202763449e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 7.964700865e-02 lcdscd = -1.416528827e-08 wcdscd = -3.122425678e-07 pcdscd = 5.957151054e-14
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 7.479338327e-01 lvoff = -1.762163339e-07 wvoff = -3.894928730e-06 pvoff = 7.704995720e-13
+ nfactor = 3.897148618e+01 lnfactor = -6.895112052e-06 wnfactor = -1.663757957e-04 pnfactor = 3.226479886e-11
+ eta0 = 8.920538562e-02 leta0 = -1.419042847e-08 weta0 = 7.142831643e-07 peta0 = -1.150317548e-13
+ etab = 5.455232265e-02 letab = -1.729337776e-08 wetab = -4.576995217e-08 petab = 1.890021661e-14
+ u0 = 8.506183898e-02 lu0 = -9.504158615e-09 wu0 = 1.060268723e-07 pu0 = -2.400614662e-14
+ ua = 6.472343722e-09 lua = -1.392789439e-15 wua = 8.242749106e-15 pua = -1.490994239e-21
+ ub = -5.052985640e-18 lub = 1.359772267e-24 wub = -5.501925139e-24 pub = 4.209306387e-31
+ uc = 1.931550608e-10 luc = -1.800861539e-17 wuc = 4.931933579e-16 puc = -1.103520864e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.603722756e+05 lvsat = -2.971981476e-02 wvsat = -1.888608824e+00 pvsat = 3.176802486e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.364558697e+00 lketa = 2.550821058e-07 wketa = 6.853085721e-06 pketa = -1.322846066e-12
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.090050787e+00 lpclm = 2.127417293e-07 wpclm = 1.380608783e-05 ppclm = -2.290297050e-12
+ pdiblc1 = -2.583725971e-01 lpdiblc1 = 1.205665408e-07 wpdiblc1 = 3.927122780e-06 ppdiblc1 = -7.475302386e-13
+ pdiblc2 = -1.070763525e-02 lpdiblc2 = 3.511295130e-09 wpdiblc2 = 1.079650739e-07 ppdiblc2 = -1.910875826e-14
+ pdiblcb = -7.100674871e-01 lpdiblcb = 1.282516707e-07 wpdiblcb = 1.109148035e-06 ppdiblcb = -2.754035238e-13
+ drout = -4.276558212e-01 ldrout = 1.782055760e-07 wdrout = 1.454870684e-05 pdrout = -2.498910068e-12
+ pscbe1 = 8.206498117e+08 lpscbe1 = -5.509145379e+00 wpscbe1 = 2.742061355e+01 ppscbe1 = 1.894360245e-7
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.677559070e-05 lalpha0 = 4.309963707e-12 walpha0 = 1.838570407e-10 palpha0 = -2.956163814e-17
+ alpha1 = 1.110374212e+01 lalpha1 = -1.648658180e-06 walpha1 = -5.571786075e-05 palpha1 = 8.958651959e-12
+ beta0 = -3.165337823e+01 lbeta0 = 7.317914033e-06 wbeta0 = 3.636407051e-04 pbeta0 = -5.846833442e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.083167237e-01 lkt1 = 7.301261631e-08 wkt1 = 7.920953037e-07 pkt1 = -1.951766773e-13
+ kt2 = -7.241605716e-02 lkt2 = 6.812207284e-09 wkt2 = 1.366762845e-09 pkt2 = 4.611276186e-16
+ at = 2.684615213e+05 lat = -4.815879108e-02 wat = -1.482757618e+00 pat = 3.090924017e-7
+ ute = -1.145774539e+01 lute = 1.842245050e-06 wute = -9.987469154e-07 pute = 1.605845215e-13
+ ua1 = -1.664587276e-08 lua1 = 3.063488002e-15 wua1 = 1.704024069e-14 pua1 = -3.206717175e-21
+ ub1 = 9.878810420e-18 lub1 = -1.646732099e-24 wub1 = -7.976112251e-24 pub1 = 1.087198166e-30
+ uc1 = 2.491233437e-10 luc1 = -7.175362263e-18 wuc1 = -1.813649820e-15 puc1 = 2.409837042e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.18 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.156258977e-01 lvth0 = 4.610520623e-08 wvth0 = -3.289744144e-09 pvth0 = 3.290098976e-13
+ k1 = 5.437593776e-01 lk1 = -2.894039739e-07 wk1 = -1.603748943e-08 pk1 = 1.603921924e-12
+ k2 = -2.747501919e-02 lk2 = 7.668108845e-08 wk2 = 5.719145794e-09 pk2 = -5.719762661e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.061689583e-01 lvoff = 9.004554036e-08 wvoff = 2.950755234e-09 pvoff = -2.951073503e-13
+ nfactor = 2.730804721e+00 lnfactor = -4.627971227e-06 wnfactor = 4.237582545e-08 pnfactor = -4.238039611e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.128149898e-02 lu0 = 1.806204949e-08 wu0 = 8.181453732e-10 pu0 = -8.182336184e-14
+ ua = -7.603977722e-10 lua = 2.438965274e-16 wua = -3.069556171e-17 pua = 3.069887253e-21
+ ub = 1.561449713e-18 lub = 9.041262229e-25 wub = 1.104602415e-25 pub = -1.104721557e-29
+ uc = 5.860591513e-11 luc = -9.364925123e-16 wuc = -4.279869903e-17 puc = 4.280331530e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.389986204e+00 la0 = -2.053741873e-06 wa0 = -1.144589624e-07 pa0 = 1.144713079e-11
+ ags = 3.837046725e-01 lags = -3.680069434e-07 wags = -2.026077567e-08 pags = 2.026296099e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.621818611e-25 lb0 = -7.622640700e-29 wb0 = -3.728541836e-30 pb0 = 3.728943997e-34
+ b1 = 2.634462122e-24 lb1 = -5.271765776e-29
+ keta = -9.255513369e-03 lketa = 4.609630834e-08 wketa = -9.360736683e-10 pketa = 9.361746332e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.607253566e-02 lpclm = 1.024456920e-06 wpclm = -1.176437843e-08 ppclm = 1.176564734e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.778937312e-03 lpdiblc2 = 2.945531555e-08 wpdiblc2 = 1.293659815e-09 ppdiblc2 = -1.293799350e-13
+ pdiblcb = -9.243755364e-01 lpdiblcb = 8.994725431e-05 wpdiblcb = 4.399683967e-06 ppdiblcb = -4.400158517e-10
+ drout = 0.56
+ pscbe1 = 8.055199410e+08 lpscbe1 = -5.085126522e+03 wpscbe1 = -1.751395166e+02 ppscbe1 = 1.751584072e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.072707742e-01 lkt1 = -5.759846956e-07 wkt1 = -1.426092497e-08 pkt1 = 1.426246316e-12
+ kt2 = -4.365554522e-02 lkt2 = -1.657970589e-07 wkt2 = -7.869767593e-09 pkt2 = 7.870616426e-13
+ at = 140000.0
+ ute = -1.762034007e+00 lute = -5.137153318e-06 wute = -1.652568725e-07 pute = 1.652746971e-11
+ ua1 = 4.312276173e-10 lua1 = -5.521357198e-15 wua1 = -1.270036222e-16 pua1 = 1.270173208e-20
+ ub1 = -6.487906259e-19 lub1 = 9.171615061e-25 wub1 = -1.286137266e-25 pub1 = 1.286275989e-29
+ uc1 = 1.485765777e-11 luc1 = 9.721600786e-17 wuc1 = 3.290266101e-18 puc1 = -3.290620990e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.19 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.179299154e-01 wvth0 = 1.315188377e-8
+ k1 = 5.292969785e-01 wk1 = 6.411538031e-8
+ k2 = -2.364303135e-02 wk2 = -2.286425249e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016691080e-01 wvoff = -1.179665900e-8
+ nfactor = 2.499530886e+00 wnfactor = -1.694119379e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.218411468e-02 wu0 = -3.270817541e-9
+ ua = -7.482095190e-10 wua = 1.227160661e-16
+ ub = 1.606631657e-18 wub = -4.416028094e-25
+ uc = 1.180652843e-11 wuc = 1.711025205e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.287354459e+00 wa0 = 4.575890716e-7
+ ags = 3.653142433e-01 wags = 8.099941968e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.047084152e-24 wb0 = 1.490612847e-29
+ b1 = 0.0
+ keta = -6.951940269e-03 wketa = 3.742276463e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.726777207e-02 wpclm = 4.703214929e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.250909254e-03 wpdiblc2 = -5.171850083e-9
+ pdiblcb = 3.570563059e+00 wpdiblcb = -1.758924998e-5
+ drout = 0.56
+ pscbe1 = 5.514006614e+08 wpscbe1 = 7.001804591e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.360544860e-01 wkt1 = 5.701295281e-8
+ kt2 = -5.194092986e-02 wkt2 = 3.146210286e-8
+ at = 140000.0
+ ute = -2.018753224e+00 wute = 6.606711901e-7
+ ua1 = 1.553085605e-10 wua1 = 5.077406641e-16
+ ub1 = -6.029572685e-19 wub1 = 5.141776104e-25
+ uc1 = 1.971583814e-11 wuc1 = -1.315397047e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.20 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.261220831e-01 lvth0 = -6.562570242e-08 wvth0 = -4.627239217e-08 pvth0 = 4.760351578e-13
+ k1 = 5.146731750e-01 lk1 = 1.171481599e-07 wk1 = 9.725702309e-08 pk1 = -2.654906080e-13
+ k2 = -2.136305342e-02 lk2 = -1.826441535e-08 wk2 = -1.900644435e-08 pk2 = -3.090407540e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.017764992e-01 lvoff = 8.602876988e-10 wvoff = -1.741041360e-08 pvoff = 4.497058676e-14
+ nfactor = 1.645326577e+00 lnfactor = 6.842847914e-06 wnfactor = 2.738429110e-06 pnfactor = -2.329409235e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.350013523e-02 lu0 = -1.054235903e-08 wu0 = -7.224255757e-09 pu0 = 3.167014752e-14
+ ua = -7.120310571e-10 lua = -2.898179157e-16 wua = -1.762999766e-17 pua = 1.124282282e-21
+ ub = 1.681817490e-18 lub = -6.022976162e-25 wub = -6.294868754e-25 pub = 1.505099045e-30
+ uc = -1.009067134e-10 luc = 9.029216596e-16 wuc = 5.270041644e-16 puc = -2.851051906e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.132572898e+00 la0 = 1.239921970e-06 wa0 = 1.075925533e-06 pa0 = -4.953361070e-12
+ ags = 2.585609582e-01 lags = 8.551777222e-07 wags = 3.059199105e-07 pags = -1.801789919e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.102384766e-24 lb0 = 2.447535939e-29 wb0 = 2.985245131e-29 pb0 = -1.197317938e-34
+ b1 = 0.0
+ keta = -1.001039642e-02 lketa = 2.450063773e-08 wketa = -1.829058468e-09 pketa = 4.463077187e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.589338897e-01 lpclm = 3.414210306e-06 wpclm = 1.042626713e-07 ppclm = -4.584614645e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 5.644443467e-03 lpdiblc2 = -1.116330436e-08 wpdiblc2 = -1.218471611e-08 ppdiblc2 = 5.617856901e-14
+ pdiblcb = 7.175821553e+00 lpdiblcb = -2.888095427e-05 wpdiblcb = -3.522592938e-05 ppdiblcb = 1.412836644e-10
+ drout = 0.56
+ pscbe1 = 3.047520763e+08 lpscbe1 = 1.975849033e+03 wpscbe1 = 1.394668907e+03 ppscbe1 = -5.563398338e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.570787832e-01 lkt1 = 1.684211460e-07 wkt1 = 1.242511916e-07 pkt1 = -5.386311418e-13
+ kt2 = -6.229710310e-02 lkt2 = 8.296108759e-08 wkt2 = 6.460144762e-08 pkt2 = -2.654721991e-13
+ at = 140000.0
+ ute = -2.359564205e+00 lute = 2.730163829e-06 wute = 1.567110738e-06 pute = -7.261293241e-12
+ ua1 = -4.790871812e-10 lua1 = 5.082008527e-15 wua1 = 2.470671323e-15 pua1 = -1.572461744e-20
+ ub1 = -1.856647873e-19 lub1 = -3.342840767e-24 wub1 = -9.084075536e-25 pub1 = 1.139602532e-29
+ uc1 = 2.750969333e-11 luc1 = -6.243490604e-17 wuc1 = -7.044317699e-17 puc1 = 4.589315736e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.21 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.849407657e-01 lvth0 = 9.954374892e-08 wvth0 = 1.493480423e-07 pvth0 = -3.085565420e-13
+ k1 = 5.392674576e-01 lk1 = 1.850575561e-08 wk1 = 2.170952134e-09 pk1 = 1.158792742e-13
+ k2 = -1.852913375e-02 lk2 = -2.963066067e-08 wk2 = -3.402362434e-08 pk2 = 2.932661985e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.297747128e+00 ldsub = -2.958945854e-06 wdsub = -2.133514529e-06 pdsub = 8.557070202e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.066412011e-01 lvoff = 2.037156588e-08 wvoff = 4.090666117e-10 pvoff = -2.649953500e-14
+ nfactor = 3.954593718e+00 lnfactor = -2.419128404e-06 wnfactor = -6.202499164e-06 pnfactor = 1.256605759e-11
+ eta0 = 2.755029890e-01 leta0 = -7.841206513e-07 weta0 = -5.653813501e-07 peta0 = 2.267623603e-12
+ etab = -2.409114178e-01 letab = 6.854891218e-07 wetab = 4.942641983e-07 petab = -1.982387927e-12
+ u0 = 3.154354951e-02 lu0 = -2.694912393e-09 wu0 = 5.497287590e-09 pu0 = -1.935324044e-14
+ ua = -7.382552809e-10 lua = -1.846381661e-16 wua = 4.229457105e-16 pua = -6.427726000e-22
+ ub = 1.498593399e-18 lub = 1.325750035e-25 wub = 8.635602547e-26 pub = -1.365993640e-30
+ uc = 1.656480202e-10 luc = -1.661723340e-16 wuc = -3.137303798e-16 puc = 5.209544339e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.129692282e+00 la0 = -2.759310497e-06 wa0 = -2.673971892e-06 pa0 = 1.008667502e-11
+ ags = 4.749010050e-01 lags = -1.251590900e-08 wags = -7.389281037e-07 pags = 2.388871869e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.063517077e-24 lb0 = -1.228711140e-29 wb0 = -1.498651722e-29 pb0 = 6.010771345e-35
+ b1 = 0.0
+ keta = -1.066710308e-02 lketa = 2.713454760e-08 wketa = 2.573665998e-08 pketa = -6.592942575e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.025958054e-01 lpclm = -4.422795344e-07 wpclm = -3.731686384e-07 ppclm = 1.456413348e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.040775976e-04 lpdiblc2 = 1.025576030e-08 wpdiblc2 = 5.269413998e-09 ppdiblc2 = -1.382621168e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.826353960e+08 lpscbe1 = 5.916130450e+01 wpscbe1 = 7.446205589e+01 ppscbe1 = -2.683311812e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.952770924e-01 lkt1 = -7.945221035e-08 wkt1 = -5.698178526e-08 pkt1 = 1.882555444e-13
+ kt2 = -4.019920264e-02 lkt2 = -5.668862200e-09 wkt2 = -7.267174950e-09 pkt2 = 2.277746618e-14
+ at = 1.624029876e+05 lat = -8.985358906e-02 wat = 7.609535152e-03 pat = -3.052021705e-8
+ ute = -1.524983364e+00 lute = -6.171613213e-07 wute = -1.204123426e-06 pute = 3.853533948e-12
+ ua1 = 1.240370863e-09 lua1 = -1.814369724e-15 wua1 = -3.515337799e-15 pua1 = 8.283984142e-21
+ ub1 = -1.494323346e-18 lub1 = 1.905908658e-24 wub1 = 3.472993146e-24 pub1 = -6.176835269e-30
+ uc1 = 3.099794454e-12 luc1 = 3.546797465e-17 wuc1 = 1.804397813e-17 puc1 = 1.040285306e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.22 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.395544222e-01 lvth0 = -1.027262686e-08 wvth0 = -1.494186265e-07 pvth0 = 2.921992927e-13
+ k1 = 4.308356169e-01 lk1 = 2.365389830e-07 wk1 = 5.829737078e-07 pk1 = -1.051990776e-12
+ k2 = 3.908106057e-03 lk2 = -7.474714835e-08 wk2 = -1.794111518e-07 pk2 = 3.216698247e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.504620890e+00 ldsub = 2.676016523e-06 wdsub = 6.847680532e-06 pdsub = -9.502191090e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -8.444723420e-02 lvoff = -2.425575203e-08 wvoff = 4.836491656e-08 pvoff = -1.229284867e-13
+ nfactor = 2.483487148e+00 lnfactor = 5.389520924e-07 wnfactor = 1.945379431e-06 pnfactor = -3.817582616e-12
+ eta0 = -2.276647030e-01 leta0 = 2.276418994e-07 weta0 = 1.116196192e-06 peta0 = -1.113668975e-12
+ etab = 7.880261914e-02 letab = 4.261261229e-08 wetab = -3.883071430e-07 petab = -2.077258298e-13
+ u0 = 3.294036187e-02 lu0 = -5.503603136e-09 wu0 = -1.632691007e-11 pu0 = -8.266541594e-15
+ ua = -3.258335162e-10 lua = -1.013930077e-15 wua = 6.515721262e-16 pua = -1.102491396e-21
+ ub = 9.565581684e-19 lub = 1.222491857e-24 wub = -1.030081871e-24 pub = 8.789240515e-31
+ uc = 1.513538305e-10 luc = -1.374297776e-16 wuc = -2.837677361e-16 puc = 4.607059694e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.398416014e+04 lvsat = 3.220442657e-02 wvsat = 5.922231393e-02 pvsat = -1.190833997e-7
+ a0 = -5.297877537e-01 la0 = 2.588334725e-06 wa0 = 7.872824655e-06 pa0 = -1.112067582e-11
+ ags = -2.734445773e-01 lags = 1.492246911e-06 wags = 7.758566726e-07 pags = -6.570361526e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.127034153e-24 lb0 = 6.193120344e-30 wb0 = 2.997303444e-29 pb0 = -3.029632359e-35
+ b1 = 0.0
+ keta = 9.607402992e-02 lketa = -1.874990283e-07 wketa = -1.255764835e-07 pketa = 2.383289247e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.242457111e+00 lpclm = -1.728903690e-06 wpclm = -3.261264820e-06 ppclm = 7.263756717e-12
+ pdiblc1 = 2.176329998e-01 lpdiblc1 = 3.465931508e-07 wpdiblc1 = -1.755111152e-07 ppdiblc1 = 3.529152932e-13
+ pdiblc2 = 3.176976609e-03 lpdiblc2 = 4.478975193e-09 wpdiblc2 = 9.421220314e-09 ppdiblc2 = -2.217460570e-14
+ pdiblcb = -5.031030115e-02 lpdiblcb = 5.089359921e-08 wpdiblcb = 6.778458428e-10 ppdiblcb = -1.363002931e-15
+ drout = 8.632358000e-01 ldrout = -6.097423013e-07 wdrout = -8.881784197e-22
+ pscbe1 = 5.779093808e+08 lpscbe1 = 4.708215096e+02 wpscbe1 = 1.705428261e+03 ppscbe1 = -3.547855193e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.347553610e-06 lalpha0 = 1.885625351e-11 walpha0 = 2.703506138e-11 palpha0 = -5.436172294e-17
+ alpha1 = 1.088945405e+00 lalpha1 = -4.804680759e-07 walpha1 = -1.337024352e-06 palpha1 = 2.688469848e-12
+ beta0 = 7.299595476e+00 lbeta0 = 1.319156957e-05 wbeta0 = 1.701667357e-05 pbeta0 = -3.421688898e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.694232834e-01 lkt1 = 6.963991258e-08 wkt1 = -5.954838544e-08 pkt1 = 1.934164281e-13
+ kt2 = -7.353752963e-02 lkt2 = 6.136737898e-08 wkt2 = 7.541524850e-08 pkt2 = -1.434791934e-13
+ at = 1.790757332e+05 lat = -1.233789125e-01 wat = -4.040650703e-02 pat = 6.602976834e-8
+ ute = -3.309734439e+00 lute = 2.971591154e-06 wute = 3.781460001e-06 pute = -6.171407408e-12
+ ua1 = -2.606269164e-09 lua1 = 5.920400189e-15 wua1 = 5.941249108e-15 pua1 = -1.073118842e-20
+ ub1 = 5.839796610e-19 lub1 = -2.273113932e-24 wub1 = 1.758326663e-25 pub1 = 4.530488623e-31
+ uc1 = -1.056356365e-10 luc1 = 2.541116569e-16 wuc1 = 6.108105077e-16 puc1 = -1.087898108e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.23 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.543335376e-01 lvth0 = 7.586745012e-08 wvth0 = 3.396081825e-07 pvth0 = -2.021021594e-13
+ k1 = 1.003286618e+00 lk1 = -3.420864745e-07 wk1 = -1.645208167e-06 pk1 = 1.200224268e-12
+ k2 = -1.865169406e-01 lk2 = 1.177318229e-07 wk2 = 5.358420685e-07 pk2 = -4.012981169e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.906612386e+00 ldsub = -7.720103144e-07 wdsub = -4.968312856e-06 pdsub = 2.441249603e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -7.604303952e-02 lvoff = -3.275059435e-08 wvoff = -1.502504314e-07 pvoff = 7.782912636e-14
+ nfactor = 3.414547571e+00 lnfactor = -4.021507483e-07 wnfactor = -4.348498945e-06 pnfactor = 2.544181532e-12
+ eta0 = -5.055270701e-01 leta0 = 5.085012900e-07 weta0 = 2.913301718e-08 peta0 = -1.488073731e-14
+ etab = 2.443880222e-01 letab = -1.247587949e-07 wetab = -1.198184333e-06 petab = 6.108866954e-13
+ u0 = 2.733751508e-02 lu0 = 1.596759531e-10 wu0 = -2.386776792e-09 pu0 = -5.870524040e-15
+ ua = -1.156606155e-09 lua = -1.741967238e-16 wua = -5.961733011e-16 pua = 1.587122137e-22
+ ub = 2.013280681e-18 lub = 1.543715351e-25 wub = 3.115756508e-25 pub = -4.772045880e-31
+ uc = -6.064487983e-11 luc = 7.685555085e-17 wuc = 3.891609163e-16 puc = -2.194808914e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.514605742e+04 lvsat = 2.092213707e-02 wvsat = -1.906577960e-01 pvsat = 1.334919171e-7
+ a0 = 2.573307362e+00 la0 = -5.482303741e-07 wa0 = -6.325869750e-06 pa0 = 3.231165706e-12
+ ags = 1.057839332e+00 lags = 1.466037740e-07 wags = 7.284138074e-07 pags = -6.090815686e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.784463315e-01 lketa = 8.998230979e-08 wketa = 3.211334837e-07 pketa = -2.131992561e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.414364367e+00 lpclm = 9.565742645e-07 wpclm = 8.107120189e-06 ppclm = -4.227247693e-12
+ pdiblc1 = -3.233753597e-01 lpdiblc1 = 8.934368265e-07 wpdiblc1 = 3.086027705e-06 ppdiblc1 = -2.943802485e-12
+ pdiblc2 = 9.495128030e-03 lpdiblc2 = -1.907323810e-09 wpdiblc2 = -1.151446740e-08 ppdiblc2 = -1.013105651e-15
+ pdiblcb = 2.562060230e-02 lpdiblcb = -2.585629497e-08 wpdiblcb = -1.355691686e-09 ppdiblcb = 6.924683333e-16
+ drout = -2.892491878e-01 ldrout = 5.551733895e-07 wdrout = -5.978030981e-07 pdrout = 6.042510023e-13
+ pscbe1 = 1.292670842e+09 lpscbe1 = -2.516493687e+02 wpscbe1 = -3.648064366e+03 ppscbe1 = 1.863380205e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.352678562e-05 lalpha0 = -1.437266833e-11 walpha0 = -7.726609104e-11 palpha0 = 5.106442172e-17
+ alpha1 = 3.721091892e-01 lalpha1 = 2.440999357e-07 walpha1 = 2.674048704e-06 palpha1 = -1.365866641e-12
+ beta0 = 3.312283359e+01 lbeta0 = -1.291019799e-05 wbeta0 = -6.407971352e-05 pbeta0 = 4.775420374e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.240128802e-01 lkt1 = 2.373971274e-08 wkt1 = 2.713191202e-07 pkt1 = -1.410198144e-13
+ kt2 = 1.032328220e-02 lkt2 = -2.339795556e-08 wkt2 = -1.302520870e-07 pkt2 = 6.440647002e-14
+ at = 4.954612963e+04 lat = 7.547797404e-03 wat = 1.027532631e-01 pat = -7.867412304e-8
+ ute = 1.078885978e+00 lute = -1.464364923e-06 wute = -6.278721734e-06 pute = 3.997283446e-12
+ ua1 = 5.529613698e-09 lua1 = -2.303236305e-15 wua1 = -9.514522320e-15 pua1 = 4.891288959e-21
+ ub1 = -1.380475416e-18 lub1 = -2.874702419e-25 wub1 = -2.768687004e-24 pub1 = 3.429328122e-30
+ uc1 = 4.034149045e-10 luc1 = -2.604295032e-16 wuc1 = -1.409192782e-15 puc1 = 9.538929368e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.24 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.680040254e-01 lvth0 = -3.327244365e-08 wvth0 = -1.342643521e-07 pvth0 = 3.994529703e-14
+ k1 = -9.599558968e-02 lk1 = 2.194114872e-07 wk1 = 1.338287641e-06 pk1 = -3.237036211e-13
+ k2 = 1.855877311e-01 lk2 = -7.233403394e-08 wk2 = -4.859201458e-07 pk2 = 1.206037176e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.000602814e-01 ldsub = 4.859400894e-08 wdsub = -6.486766524e-07 pdsub = 2.348399052e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.399062768e-01 lvoff = -1.301468342e-10 wvoff = 1.834511416e-08 pvoff = -8.287117955e-15
+ nfactor = 2.100585880e+00 lnfactor = 2.690024878e-07 wnfactor = 1.253257892e-06 pnfactor = -3.171174356e-13
+ eta0 = 0.49
+ etab = 2.143669139e-03 letab = -1.023770813e-09 wetab = -8.006802879e-09 petab = 2.960675575e-15
+ u0 = 3.841614930e-02 lu0 = -5.499135301e-09 wu0 = -2.132978318e-08 pu0 = 3.805298420e-15
+ ua = -8.244069547e-10 lua = -3.438794247e-16 wua = -7.543233911e-16 pua = 2.394930655e-22
+ ub = 2.052005131e-18 lub = 1.345916279e-25 wub = -3.208321031e-25 pub = -1.541795610e-31
+ uc = 1.741587971e-10 luc = -4.307888005e-17 wuc = -2.802302278e-16 puc = 1.224347335e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.042416423e+05 lvsat = 6.060519664e-03 wvsat = -4.539936912e-02 pvsat = 5.929594623e-8
+ a0 = 1.5
+ ags = 2.727358896e+00 lags = -7.061634462e-07 wags = -9.480701297e-07 pags = 2.472429557e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.763841729e-02 lketa = -1.017503471e-08 wketa = -1.407424350e-07 pketa = 2.272049684e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.358960122e-01 lpclm = 6.256576657e-08 wpclm = 4.227082817e-07 ppclm = -3.021576722e-13
+ pdiblc1 = 1.872845312e+00 lpdiblc1 = -2.283619457e-07 wpdiblc1 = -2.930628606e-06 ppdiblc1 = 1.294213259e-13
+ pdiblc2 = 9.203791952e-03 lpdiblc2 = -1.758513420e-09 wpdiblc2 = -2.794247220e-08 ppdiblc2 = 7.378089205e-15
+ pdiblcb = -3.266701514e-01 lpdiblcb = 1.540888900e-07 wpdiblcb = 1.475749867e-06 ppdiblcb = -7.537923717e-13
+ drout = 5.865718156e-01 ldrout = 1.078162825e-07 wdrout = 1.195606196e-06 pdrout = -3.117973575e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.592623138e-05 lalpha0 = 5.779380403e-12 walpha0 = 5.524643575e-11 palpha0 = -1.662112180e-17
+ alpha1 = 0.85
+ beta0 = -4.625052572e+00 lbeta0 = 6.370893794e-06 wbeta0 = 6.213664633e-05 pbeta0 = -1.671534584e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.405920253e-01 lkt1 = -1.887049208e-08 wkt1 = -2.107395881e-07 pkt1 = 1.052090250e-13
+ kt2 = -3.085713183e-02 lkt2 = -2.363576601e-09 wkt2 = -7.730641724e-08 pkt2 = 3.736256315e-14
+ at = 9.628588818e+04 lat = -1.632621690e-02 wat = -7.160444954e-02 pat = 1.038535556e-8
+ ute = -2.438414063e+00 lute = 3.322226955e-07 wute = 4.942141822e-07 pute = 5.377626013e-13
+ ua1 = 1.384509975e-09 lua1 = -1.859753549e-16 wua1 = -5.053915635e-15 pua1 = 2.612873513e-21
+ ub1 = -3.941920592e-18 lub1 = 1.020880094e-24 wub1 = 1.233486838e-23 pub1 = -4.285356519e-30
+ uc1 = -3.437286223e-10 luc1 = 1.212009503e-16 wuc1 = 1.148336553e-15 puc1 = -3.524572421e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.25 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 7.730160506e-01 lvth0 = -6.065810965e-08 wvth0 = -5.209818835e-07 pvth0 = 1.407958152e-13
+ k1 = 4.371245774e-01 lk1 = 8.038121129e-08 wk1 = -2.185173437e-08 pk1 = 3.100168605e-14
+ k2 = 5.507251898e-04 lk2 = -2.407897333e-08 wk2 = 1.231549536e-07 pk2 = -3.823454132e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 9.846145802e-01 ldsub = -1.299281684e-07 wdsub = -2.837501014e-07 pdsub = 1.396721697e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -7.794471313e-03 lcdscd = 3.440933396e-09 wcdscd = 6.454645644e-08 pcdscd = -1.683281219e-14
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.649240481e-01 lvoff = 3.247273768e-08 wvoff = 6.382217716e-07 pvoff = -1.699422719e-13
+ nfactor = -9.830844703e-01 lnfactor = 1.073180544e-06 wnfactor = 1.681925887e-05 pnfactor = -4.376512567e-12
+ eta0 = 1.577656670e+00 leta0 = -2.836456324e-07 weta0 = 7.112806273e-07 peta0 = -1.854920297e-13
+ etab = -4.029506008e-02 letab = 1.004365563e-08 wetab = 5.130479682e-07 petab = -1.329231140e-13
+ u0 = -2.933691754e-02 lu0 = 1.216991599e-08 wu0 = 1.826920525e-08 pu0 = -6.521563375e-15
+ ua = -7.727338474e-09 lua = 1.456308474e-15 wua = 9.228952702e-15 pua = -2.364005574e-21
+ ub = 7.940176805e-18 lub = -1.400961110e-24 wub = -1.411045937e-23 pub = 3.441962174e-30
+ uc = -2.734310462e-10 luc = 7.364628480e-17 wuc = 1.121591051e-15 puc = -2.431406306e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.483384794e+05 lvsat = -5.439318103e-03 wvsat = 1.568731938e-01 pvsat = 6.546093629e-9
+ a0 = 1.5
+ ags = -3.334127560e+00 lags = 8.745873606e-07 wags = -6.588169051e-12 pags = 1.256930421e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.387875616e-02 lketa = -9.194567721e-09 wketa = -7.030020982e-08 pketa = 4.350150714e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.294973822e-01 lpclm = 1.207723970e-08 wpclm = -8.179378332e-08 ppclm = -1.705905967e-13
+ pdiblc1 = 2.619177152e+00 lpdiblc1 = -4.229948409e-07 wpdiblc1 = -8.713837152e-06 ppdiblc1 = 1.637601150e-12
+ pdiblc2 = -1.965367562e-02 lpdiblc2 = 5.767110119e-09 wpdiblc2 = 1.839232551e-08 ppdiblc2 = -4.705377350e-15
+ pdiblcb = 1.285093666e+00 lpdiblcb = -2.662365489e-07 wpdiblcb = -5.326361177e-06 ppdiblcb = 1.020102959e-12
+ drout = 3.561772454e-01 ldrout = 1.678999609e-07 wdrout = 5.776671875e-06 pdrout = -1.506475152e-12
+ pscbe1 = 7.823053059e+08 lpscbe1 = 4.614528506e+00 wpscbe1 = 1.188003750e+02 ppscbe1 = -3.098147460e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.184899916e-05 lalpha0 = -1.464010867e-12 walpha0 = 1.051022245e-12 palpha0 = -2.487716688e-18
+ alpha1 = 2.040839624e+00 lalpha1 = -3.105543021e-07 walpha1 = -3.443827214e-06 palpha1 = 8.981019240e-13
+ beta0 = 7.330784214e+00 lbeta0 = 3.252978942e-06 wbeta0 = 7.255437756e-05 pbeta0 = -1.943214430e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.361396470e-01 lkt1 = 6.046990006e-09 wkt1 = 2.963136104e-07 pkt1 = -2.702335043e-14
+ kt2 = -2.296425315e-02 lkt2 = -4.421928863e-09 wkt2 = 1.096797691e-07 pkt2 = -1.140081644e-14
+ at = 1.298124945e+05 lat = -2.506948646e-02 wat = -7.277514404e-01 pat = 1.814993047e-7
+ ute = 2.688182574e+00 lute = -1.004721935e-06 wute = -3.999067216e-07 pute = 7.709368153e-13
+ ua1 = 6.015080865e-09 lua1 = -1.393563415e-15 wua1 = 8.524450261e-15 pua1 = -9.281742155e-22
+ ub1 = -2.525137353e-18 lub1 = 6.514028599e-25 wub1 = -1.383568890e-23 pub1 = 2.539558431e-30
+ uc1 = 3.711290816e-10 luc1 = -6.522393088e-17 wuc1 = -1.686458139e-15 puc1 = 3.868175264e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.26 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.149419683e-01 lvth0 = -1.142118778e-08 wvth0 = 4.538638783e-07 pvth0 = -4.519110833e-14
+ k1 = 6.685934923e-01 lk1 = 3.622018288e-08 wk1 = 6.896679366e-07 pk1 = -1.047463059e-13
+ k2 = -9.081029267e-02 lk2 = -6.648570177e-09 wk2 = -9.400709982e-08 pk2 = 3.196938201e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.380909432e-01 ldsub = -6.580509818e-09 wdsub = 3.486673228e-07 pdsub = 1.901577900e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 3.572544955e-02 lcdscd = -4.862058226e-09 wcdscd = -9.738132631e-08 pcdscd = 1.406074177e-14
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 1.451800107e-01 lvoff = -4.576937528e-08 wvoff = -9.462980199e-07 pvoff = 1.323619210e-13
+ nfactor = 1.284791319e+01 lnfactor = -1.565580175e-06 wnfactor = -3.858105295e-05 pnfactor = 6.193091324e-12
+ eta0 = 5.743312101e-01 leta0 = -9.222518117e-08 weta0 = -1.658919380e-06 peta0 = 2.667089490e-13
+ etab = 1.845252169e-01 letab = -3.284890573e-08 wetab = -6.815885125e-07 petab = 9.499680166e-14
+ u0 = 2.268845522e-01 lu0 = -3.671355334e-08 wu0 = -5.877601969e-07 pu0 = 1.091003621e-13
+ ua = 2.167070205e-08 lua = -4.152426084e-15 wua = -6.610658633e-14 pua = 1.200896058e-20
+ ub = -1.779112800e-17 lub = 3.508211608e-24 wub = 5.681220109e-23 pub = -1.008908852e-29
+ uc = 6.326668275e-10 luc = -9.922450413e-17 wuc = -1.656868318e-15 puc = 2.869505187e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.186456878e+05 lvsat = 6.457612321e-02 wvsat = 9.439076799e-01 pvsat = -1.436090678e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.981917596e-01 lketa = -1.397519084e-07 wketa = -3.237749247e-06 pketa = 6.086550827e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.125584191e+00 lpclm = -4.832197783e-07 wpclm = -6.816511825e-06 ppclm = 1.114299320e-12
+ pdiblc1 = 8.154212105e-01 lpdiblc1 = -7.886345980e-08 wpdiblc1 = -1.325803508e-06 ppdiblc1 = 2.280677630e-13
+ pdiblc2 = 1.563707289e-02 lpdiblc2 = -9.658706263e-10 wpdiblc2 = -2.091144689e-08 ppdiblc2 = 2.793232172e-15
+ pdiblcb = -1.032864742e+00 lpdiblcb = 1.759974640e-07 wpdiblcb = 2.688250257e-06 ppdiblcb = -5.089726980e-13
+ drout = 5.500528586e+00 ldrout = -8.135702539e-07 wdrout = -1.445156816e-05 pdrout = 2.352789852e-12
+ pscbe1 = 8.766256060e+08 lpscbe1 = -1.338046427e+01 wpscbe1 = -2.464091656e+02 ppscbe1 = 3.869539281e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.639295687e-05 lalpha0 = -4.238794384e-12 walpha0 = -7.623987860e-11 palpha0 = 1.225830512e-17
+ alpha1 = -1.928625788e+00 lalpha1 = 4.467641260e-07 walpha1 = 8.035596834e-06 palpha1 = -1.292011473e-12
+ beta0 = 8.076986596e+01 lbeta0 = -1.075816971e-05 wbeta0 = -1.863261607e-04 pbeta0 = 2.995863807e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.289936741e-01 lkt1 = 8.099803842e-08 wkt1 = 1.382438739e-06 pkt1 = -2.342408193e-13
+ kt2 = -1.346858683e-01 lkt2 = 1.689299121e-08 wkt2 = 3.059864447e-07 pkt2 = -4.885338186e-14
+ at = -3.104658499e+05 lat = 5.892945775e-02 wat = 1.349315715e+00 pat = -2.147760296e-7
+ ute = -2.661733750e+01 lute = 4.586361017e-06 wute = 7.316094682e-05 pute = -1.326344419e-11
+ ua1 = -3.216063602e-08 lua1 = 5.889828907e-15 wua1 = 9.293740757e-14 pua1 = -1.703298469e-20
+ ub1 = 1.915179126e-17 lub1 = -3.484251643e-24 wub1 = -5.333890397e-23 pub1 = 1.007621882e-29
+ uc1 = -5.103039945e-10 luc1 = 1.029411600e-16 wuc1 = 1.901417078e-15 puc1 = -2.976988347e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.27 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.037705701e-01 lvth0 = 3.743443722e-07 wvth0 = 3.099505687e-08 pvth0 = -6.202354501e-13
+ k1 = 5.345769059e-01 lk1 = 3.379922632e-07 wk1 = 1.051759441e-08 pk1 = -2.104653309e-13
+ k2 = -2.169276183e-02 lk2 = -1.972361156e-07 wk2 = -1.100274930e-08 pk2 = 2.201736616e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.079585345e-01 lvoff = 4.422912971e-08 wvoff = 8.126087911e-09 pvoff = -1.626094062e-13
+ nfactor = 3.264920145e+00 lnfactor = -1.648829025e-05 wnfactor = -1.502249661e-06 pnfactor = 3.006119649e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.143810506e-02 lu0 = -7.704253888e-09 wu0 = 3.652512495e-10 pu0 = -7.308964590e-15
+ ua = -8.534025596e-10 lua = 2.954131897e-15 wua = 2.382679590e-16 pua = -4.767929139e-21
+ ub = 1.727672372e-18 lub = -5.477800018e-24 wub = -3.702443845e-25 pub = 7.408881147e-30
+ uc = 4.962252348e-11 luc = 4.272198059e-16 wuc = -1.681934124e-17 puc = 3.365682383e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.323342844e+00 la0 = 2.446141610e-06 wa0 = 7.826910202e-08 pa0 = -1.566226251e-12
+ ags = 3.723302380e-01 lags = 4.200816687e-07 wags = 1.263331569e-08 pags = -2.528025767e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.271091167e-25 lb0 = 5.271659707e-29
+ b1 = 7.618685315e-24 lb1 = -1.524558814e-28 wb1 = -1.441403454e-29 pb1 = 2.884361607e-34
+ keta = -1.574673177e-02 lketa = 2.018854536e-07 wketa = 1.783608855e-08 pketa = -3.569141510e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.075926543e-01 lpclm = 3.824534545e-06 wpclm = 3.458669416e-07 ppclm = -6.921069353e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.941906546e-03 lpdiblc2 = -9.592555392e-09 wpdiblc2 = 8.223638722e-10 ppdiblc2 = -1.645614746e-14
+ pdiblcb = 5.969894081e-01 lpdiblcb = -6.220564959e-05 wpdiblcb = 1.942890293e-22 ppdiblcb = 9.769962617e-27
+ drout = 0.56
+ pscbe1 = 8.872089763e+08 lpscbe1 = -1.874874501e+03 wpscbe1 = -4.113786519e+02 ppscbe1 = 8.232010169e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.853100699e-01 lkt1 = -6.209332904e-07 wkt1 = -7.776978851e-08 pkt1 = 1.556234595e-12
+ kt2 = -4.591286303e-02 lkt2 = 9.707634562e-08 wkt2 = -1.341757989e-09 pkt2 = 2.684963198e-14
+ at = 140000.0
+ ute = -1.652906658e+00 lute = -2.749348768e-06 wute = -4.808457460e-07 pute = 9.622101323e-12
+ ua1 = 6.638467717e-10 lua1 = -6.662926814e-15 wua1 = -7.997223987e-16 pua1 = 1.600307378e-20
+ ub1 = -1.028574077e-18 lub1 = 1.207478996e-23 wub1 = 9.696941880e-25 pub1 = -1.940434288e-29
+ uc1 = 1.316378282e-11 luc1 = 4.009259381e-17 wuc1 = 8.188837255e-18 puc1 = -1.638650699e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.28 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.5224777
+ k1 = 0.55146741
+ k2 = -0.031549252
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10574827
+ nfactor = 2.44095
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0310531
+ ua = -7.0577558e-10
+ ub = 1.45393e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.445584
+ ags = 0.393323
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.29 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.101215713e-01 lvth0 = 9.898230280e-8
+ k1 = 5.483036418e-01 lk1 = 2.534426967e-8
+ k2 = -2.793528414e-02 lk2 = -2.895072312e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.077968391e-01 lvoff = 1.641064876e-8
+ nfactor = 2.592246875e+00 lnfactor = -1.212006887e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.100206275e-02 lu0 = 4.088485026e-10
+ ua = -7.181273269e-10 lua = 9.894720127e-17
+ ub = 1.464147477e-18 lub = -8.185002439e-26
+ uc = 8.132584406e-11 luc = -8.294242903e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.504616754e+00 la0 = -4.728987572e-7
+ ags = 3.643448806e-01 lags = 2.321375129e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.220282334e-24 lb0 = -1.692664930e-29
+ b1 = 0.0
+ keta = -1.064286581e-02 lketa = 3.993349433e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.228809427e-01 lpclm = 3.255679101e-06 wpclm = -1.110223025e-22 ppclm = 1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.431095396e-03 lpdiblc2 = 8.262660361e-9
+ pdiblcb = -5.004938362e+00 lpdiblcb = 1.997346706e-05 ppdiblcb = 1.421085472e-26
+ drout = 0.56
+ pscbe1 = 7.870140753e+08 lpscbe1 = 5.208376498e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141140138e-01 lkt1 = -1.783189933e-8
+ kt2 = -3.995859458e-02 lkt2 = -8.836437064e-9
+ at = 140000.0
+ ute = -1.817673614e+00 lute = 2.192841674e-7
+ ua1 = 3.752452592e-10 lua1 = -3.554005973e-16
+ ub1 = -4.997826689e-19 lub1 = 5.977862313e-25
+ uc1 = 3.151175570e-12 luc1 = 9.625885770e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.30 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.365837650e-01 lvth0 = -7.151893317e-9
+ k1 = 5.400181503e-01 lk1 = 5.857560310e-8
+ k2 = -3.029414909e-02 lk2 = -1.948982062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.064997501e-01 lvoff = 1.120830236e-8
+ nfactor = 1.809834034e+00 lnfactor = 1.926083583e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.344445436e-02 lu0 = -9.387061600e-9
+ ua = -5.920050542e-10 lua = -4.069022443e-16
+ ub = 1.528454414e-18 lub = -3.397713864e-25
+ uc = 5.716331865e-11 luc = 1.396828961e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205060620e+00 la0 = 7.285567913e-7
+ ags = 2.193873541e-01 lags = 8.135311311e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.118664669e-24 lb0 = 8.497510593e-30
+ b1 = 0.0
+ keta = -1.767633807e-03 lketa = 4.336838064e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.735579725e-01 lpclm = 6.133304993e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.126186139e-03 lpdiblc2 = 5.474800142e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.083836002e+08 lpscbe1 = -3.362482644e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.149808009e-01 lkt1 = -1.435540156e-8
+ kt2 = -4.271211613e-02 lkt2 = 2.207348643e-9
+ at = 1.650342857e+05 lat = -1.004071626e-1
+ ute = -1.941356718e+00 lute = 7.153506284e-7
+ ua1 = 2.480362285e-11 lua1 = 1.050145812e-15
+ ub1 = -2.933984465e-19 lub1 = -2.299767186e-25
+ uc1 = 9.339214374e-12 luc1 = 7.143995830e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.31 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.878870156e-01 lvth0 = 9.076684872e-8
+ k1 = 6.324218602e-01 lk1 = -1.272284831e-7
+ k2 = -5.813040379e-02 lk2 = 3.648293062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.772314921e-02 lvoff = -6.676314387e-8
+ nfactor = 3.156179117e+00 lnfactor = -7.811282609e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 3.293471619e-02 lu0 = -8.362087220e-9
+ ua = -1.005266535e-10 lua = -1.395160132e-15
+ ub = 6.003665738e-19 lub = 1.526414650e-24
+ uc = 5.322989950e-11 luc = 2.187755377e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.446262019e+04 lvsat = -8.973374201e-3
+ a0 = 2.192553109e+00 la0 = -1.257079281e-6
+ ags = -5.161411334e-03 lags = 1.265050645e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.237329338e-24 lb0 = -4.283033172e-30
+ b1 = 0.0
+ keta = 5.265098834e-02 lketa = -1.050873655e-07 wketa = 1.647987302e-23 pketa = -5.464378949e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.147456642e-01 lpclm = 7.828278159e-7
+ pdiblc1 = 1.569430821e-01 lpdiblc1 = 4.686275877e-7
+ pdiblc2 = 6.434736582e-03 lpdiblc2 = -3.188772769e-9
+ pdiblcb = -5.007590911e-02 lpdiblcb = 5.042228697e-8
+ drout = 8.632358000e-01 ldrout = -6.097423013e-7
+ pscbe1 = 1.167628731e+09 lpscbe1 = -7.559899069e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 8.893632000e-10 lalpha0 = 5.853526093e-14
+ alpha1 = 6.266162940e-01 lalpha1 = 4.491768287e-7
+ beta0 = 1.318378417e+01 lbeta0 = 1.359725332e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.900144956e-01 lkt1 = 1.365213013e-7
+ kt2 = -4.745972127e-02 lkt2 = 1.175376658e-8
+ at = 1.651035834e+05 lat = -1.005465055e-1
+ ute = -2.002144911e+00 lute = 8.375826746e-7
+ ua1 = -5.518470310e-10 lua1 = 2.209666873e-15
+ ub1 = 6.447807678e-19 lub1 = -2.116454348e-24
+ uc1 = 1.055762826e-10 luc1 = -1.220721912e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.32 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.717665141e-01 lvth0 = 5.982625921e-9
+ k1 = 4.343907494e-01 lk1 = 7.293859126e-8
+ k2 = -1.228327853e-03 lk2 = -2.103289110e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.886214874e-01 ldsub = 7.214840124e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.279980756e-01 lvoff = -5.838092139e-9
+ nfactor = 1.910881874e+00 lnfactor = 4.776007576e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 6.938893904e-23 peta0 = 1.786765180e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.651219250e-02 lu0 = -1.870290187e-9
+ ua = -1.362756681e-09 lua = -1.193156915e-16
+ ub = 2.121020299e-18 lub = -1.064084691e-26
+ uc = 7.392291647e-11 luc = 9.613419190e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.218575020e+03 lvsat = 6.708225324e-2
+ a0 = 3.858874119e-01 la0 = 5.690731124e-7
+ ags = 1.309717248e+00 lags = -6.401029598e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.740171369e-02 lketa = 1.626022499e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.388993454e+00 lpclm = -5.051640103e-7
+ pdiblc1 = 7.437409158e-01 lpdiblc1 = -1.244994474e-07 wpdiblc1 = 8.881784197e-22
+ pdiblc2 = 5.513544990e-03 lpdiblc2 = -2.257645204e-9
+ pdiblcb = 2.515181822e-02 lpdiblcb = -2.561684662e-08 wpdiblcb = 1.214306433e-23 ppdiblcb = 2.168404345e-31
+ drout = -4.959632800e-01 ldrout = 7.641170999e-7
+ pscbe1 = 3.120813611e+07 lpscbe1 = 3.926881210e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.191024846e-06 lalpha0 = 3.284877457e-12 walpha0 = -1.482307658e-27 palpha0 = 7.411538288e-34
+ alpha1 = 1.296767412e+00 lalpha1 = -2.282025393e-7
+ beta0 = 1.096473529e+01 lbeta0 = 3.602708867e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.301935511e-01 lkt1 = -2.502347200e-8
+ kt2 = -3.471653443e-02 lkt2 = -1.126868269e-9
+ at = 8.507713903e+04 lat = -1.965689587e-2
+ ute = -1.092230678e+00 lute = -8.214589253e-8
+ ua1 = 2.239590862e-09 lua1 = -6.118794686e-16
+ ub1 = -2.337858579e-18 lub1 = 8.983557464e-25
+ uc1 = -8.386929930e-11 luc1 = 6.941675076e-17 wuc1 = 2.584939414e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.33 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.215768093e-01 lvth0 = -1.945977550e-8
+ k1 = 3.667703539e-01 lk1 = 1.074781426e-7
+ k2 = 1.756159980e-02 lk2 = -3.063052309e-08 pk2 = 1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 7.575464332e-02 ldsub = 1.297992051e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.335627272e-01 lvoff = -2.995746010e-9
+ nfactor = 2.533949421e+00 lnfactor = 1.593465777e-7
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 3.104053217e-02 lu0 = -4.183302695e-9
+ ua = -1.085244136e-09 lua = -2.610652142e-16
+ ub = 1.941064728e-18 lub = 8.127793964e-26
+ uc = 7.725809959e-11 luc = -7.422229282e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.854301274e+04 lvsat = 2.656444100e-2
+ a0 = 1.5
+ ags = 2.399526108e+00 lags = -6.206694043e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.102885254e-02 lketa = -2.318523268e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.820641385e-01 lpclm = -4.191721304e-8
+ pdiblc1 = 8.594644286e-01 lpdiblc1 = -1.836093976e-7
+ pdiblc2 = -4.584242403e-04 lpdiblc2 = 7.927530709e-10 ppdiblc2 = 4.336808690e-31
+ pdiblcb = 1.836288000e-01 lpdiblcb = -1.065646702e-07 wpdiblcb = -1.110223025e-22
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.177411360e-06 lalpha0 = 3.196940107e-14
+ alpha1 = 0.85
+ beta0 = 1.686115330e+01 lbeta0 = 5.909010965e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.134635824e-01 lkt1 = 1.750969425e-8
+ kt2 = -5.758888667e-02 lkt2 = 1.055600904e-8
+ at = 7.152581445e+04 lat = -1.273506899e-2
+ ute = -2.267519941e+00 lute = 5.181754085e-7
+ ua1 = -3.630814747e-10 lua1 = 7.175291234e-16
+ ub1 = 3.233485706e-19 lub1 = -4.609516086e-25 pub1 = -1.925929944e-46
+ uc1 = 5.335421127e-11 luc1 = -6.750973096e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.34 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.826818720e-01 lvth0 = -9.316520387e-09 wvth0 = 2.945161824e-08 pvth0 = -7.680569715e-15
+ k1 = 4.295684749e-01 lk1 = 9.110127180e-8
+ k2 = 6.613024587e-03 lk2 = -2.777528795e-08 wk2 = 1.056231960e-07 pk2 = -2.754505078e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.864712740e-01 ldsub = -8.162434218e-08 wdsub = 7.366632614e-11 pdsub = -1.921114653e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.452502183e-02 lcdscd = -2.379677943e-09 wcdscd = -1.387778781e-23
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.756724704e-01 lvoff = 7.985885496e-09 wvoff = 3.801122780e-07 pvoff = -9.912796053e-14
+ nfactor = 2.349537676e+00 lnfactor = 2.074385790e-07 wnfactor = 7.181542241e-06 pnfactor = -1.872845675e-12
+ eta0 = 1.823610105e+00 leta0 = -3.477868449e-07 weta0 = 1.819289785e-14 peta0 = -4.744453275e-21
+ etab = 1.740475113e-01 letab = -4.555214553e-08 wetab = -1.068161729e-07 petab = 2.785616247e-14
+ u0 = -1.260304720e-02 lu0 = 7.198331796e-09 wu0 = -3.012400987e-08 pu0 = 7.855920038e-15
+ ua = -4.266324707e-09 lua = 5.685160635e-16 wua = -7.800637625e-16 pua = 2.034297084e-22
+ ub = 1.928304229e-18 lub = 8.460569905e-26 wub = 3.275467315e-24 pub = -8.541960192e-31
+ uc = 2.314608982e-10 luc = -4.095615398e-17 wuc = -3.385221194e-16 puc = 8.828182942e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.036146612e+05 lvsat = -2.952323392e-02 wvsat = -2.921749652e-01 pvsat = 7.619514047e-8
+ a0 = 1.5
+ ags = -3.334129838e+00 lags = 8.745877952e-07 wags = -5.551115123e-22 pags = -3.330669074e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.461768944e-01 lketa = -1.006885012e-07 wketa = -1.031283829e-06 pketa = 2.689443847e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.541814529e-02 lpclm = 9.042706182e-08 wpclm = 1.522984188e-06 ppclm = -3.971729544e-13
+ pdiblc1 = -3.939770822e-01 lpdiblc1 = 1.432706002e-7
+ pdiblc2 = -1.329380080e-02 lpdiblc2 = 4.140039583e-09 wpdiblc2 = 6.938893904e-24 ppdiblc2 = -1.734723476e-30
+ pdiblcb = -5.567066175e-01 lpdiblcb = 8.650444195e-8
+ drout = 2.353690284e+00 ldrout = -3.530234743e-7
+ pscbe1 = 8.233852396e+08 lpscbe1 = -6.098543103e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.221243171e-05 lalpha0 = -2.324237417e-12
+ alpha1 = 0.85
+ beta0 = 3.040830297e+01 lbeta0 = -2.942005877e-06 wbeta0 = 5.815762590e-06 pbeta0 = -1.516669463e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.821126062e-01 lkt1 = -1.674480144e-08 wkt1 = -1.491221177e-07 pkt1 = 3.888896058e-14
+ kt2 = 1.496186997e-02 lkt2 = -8.364212580e-9
+ at = -1.991836980e+05 lat = 5.786218192e-02 wat = 2.236831765e-01 pat = -5.833344087e-8
+ ute = 2.549898990e+00 lute = -7.381400046e-07 pute = 4.440892099e-28
+ ua1 = 8.962747083e-09 lua1 = -1.714516403e-15
+ ub1 = -7.309374636e-18 lub1 = 1.529555746e-24
+ uc1 = -2.120305980e-10 luc1 = 6.853354557e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.35 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 9.438398519e-01 lvth0 = -7.822040675e-08 wvth0 = -7.864796361e-07 pvth0 = 1.479876906e-13
+ k1 = 0.90707349
+ k2 = -5.494816598e-02 lk2 = -1.603027465e-08 wk2 = -1.977179316e-07 pk2 = 3.032818958e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587159132e-01 ldsub = -1.460792414e-11 wdsub = -1.718880943e-10 pdsub = 2.763719913e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.338146533e-01 wvoff = -1.394644233e-7
+ nfactor = -5.293063660e+00 lnfactor = 1.665539917e-06 wnfactor = 1.388141850e-05 pnfactor = -3.151088267e-12
+ eta0 = 6.941612174e-04 leta0 = -3.607624990e-15 weta0 = -4.245009617e-14 peta0 = 6.825381162e-21
+ etab = -6.471290892e-02 wetab = 3.919119906e-8
+ u0 = 9.783655146e-03 lu0 = 2.927262402e-09 wu0 = 4.008083455e-08 pu0 = -5.538181410e-15
+ ua = -1.288698684e-09 lua = 4.267051525e-19 wua = 2.904393431e-16 pua = -8.072971326e-25
+ ub = 2.076034198e-18 lub = 5.642088919e-26 wub = -6.422810181e-25 pub = -1.067444857e-31
+ uc = 1.679025167e-11 wuc = 1.242048597e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.725145711e+04 lvsat = 4.314068933e-02 wvsat = 5.350051796e-01 pvsat = -8.161925064e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.253471759e+00 lketa = 2.045020667e-07 wketa = 2.406328935e-06 pketa = -3.869040041e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.932621135e+00 lpclm = -2.831394203e-07 wpclm = -3.366543787e-06 ppclm = 5.356805298e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 2.103262180e+01 lbeta0 = -1.153257169e-06 wbeta0 = -1.357011271e-05 pbeta0 = 2.181884142e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.698800600e-01 wkt1 = 5.471338693e-8
+ kt2 = -0.028878939
+ at = 3.365905563e+05 lat = -4.435604496e-02 wat = -5.219274119e-01 pat = 8.391862085e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.36 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.201533243e-01 lvth0 = 4.651258432e-8
+ k1 = 5.401360879e-01 lk1 = 2.267486609e-7
+ k2 = -2.750837745e-02 lk2 = -8.086107591e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.036634077e-01 lvoff = -4.171973431e-8
+ nfactor = 2.470890729e+00 lnfactor = -5.991375219e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.163116234e-02 lu0 = -1.156748184e-8
+ ua = -7.274635940e-10 lua = 4.339942073e-16
+ ub = 1.531975917e-18 lub = -1.561760146e-24
+ uc = 4.073248872e-11 luc = 6.051163890e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.364712778e+00 la0 = 1.618296714e-6
+ ags = 3.790077061e-01 lags = 2.864602824e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.271091167e-25 lb0 = 5.271659707e-29
+ b1 = 0.0
+ keta = -6.319284829e-03 lketa = 1.323483028e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.521885355e-02 lpclm = 1.663325838e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.376575378e-03 lpdiblc2 = -1.829062036e-8
+ pdiblcb = 5.969894081e-01 lpdiblcb = -6.220564959e-05 wpdiblcb = -2.775557562e-22 ppdiblcb = -3.907985047e-26
+ drout = 0.56
+ pscbe1 = 6.697705843e+08 lpscbe1 = 2.476238630e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.264160867e-01 lkt1 = 2.016304145e-7
+ kt2 = -4.662206293e-02 lkt2 = 1.112679931e-7
+ at = 140000.0
+ ute = -1.907062593e+00 lute = 2.336511254e-6
+ ua1 = 2.411453223e-10 lua1 = 1.795661433e-15
+ ub1 = -5.160323004e-19 lub1 = 1.818426157e-24
+ uc1 = 1.749207647e-11 luc1 = -4.651996409e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.37 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.5224777
+ k1 = 0.55146741
+ k2 = -0.031549252
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10574827
+ nfactor = 2.44095
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0310531
+ ua = -7.0577558e-10
+ ub = 1.45393e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.445584
+ ags = 0.393323
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.38 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.101215713e-01 lvth0 = 9.898230280e-8
+ k1 = 5.483036418e-01 lk1 = 2.534426967e-8
+ k2 = -2.793528414e-02 lk2 = -2.895072312e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.077968391e-01 lvoff = 1.641064876e-8
+ nfactor = 2.592246875e+00 lnfactor = -1.212006887e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.100206275e-02 lu0 = 4.088485026e-10
+ ua = -7.181273269e-10 lua = 9.894720127e-17
+ ub = 1.464147477e-18 lub = -8.185002439e-26
+ uc = 8.132584406e-11 luc = -8.294242903e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.504616754e+00 la0 = -4.728987572e-7
+ ags = 3.643448806e-01 lags = 2.321375129e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.220282334e-24 lb0 = -1.692664930e-29
+ b1 = 0.0
+ keta = -1.064286581e-02 lketa = 3.993349433e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.228809427e-01 lpclm = 3.255679101e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.431095396e-03 lpdiblc2 = 8.262660361e-9
+ pdiblcb = -5.004938362e+00 lpdiblcb = 1.997346706e-5
+ drout = 0.56
+ pscbe1 = 7.870140753e+08 lpscbe1 = 5.208376498e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141140138e-01 lkt1 = -1.783189933e-8
+ kt2 = -3.995859458e-02 lkt2 = -8.836437064e-9
+ at = 140000.0
+ ute = -1.817673614e+00 lute = 2.192841674e-7
+ ua1 = 3.752452592e-10 lua1 = -3.554005973e-16
+ ub1 = -4.997826689e-19 lub1 = 5.977862313e-25
+ uc1 = 3.151175570e-12 luc1 = 9.625885770e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.39 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.365837650e-01 lvth0 = -7.151893317e-9
+ k1 = 5.400181503e-01 lk1 = 5.857560310e-8
+ k2 = -3.029414909e-02 lk2 = -1.948982062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.064997501e-01 lvoff = 1.120830236e-8
+ nfactor = 1.809834034e+00 lnfactor = 1.926083583e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.344445436e-02 lu0 = -9.387061600e-9
+ ua = -5.920050542e-10 lua = -4.069022443e-16
+ ub = 1.528454414e-18 lub = -3.397713864e-25
+ uc = 5.716331865e-11 luc = 1.396828961e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205060620e+00 la0 = 7.285567913e-7
+ ags = 2.193873541e-01 lags = 8.135311311e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.118664669e-24 lb0 = 8.497510593e-30
+ b1 = 0.0
+ keta = -1.767633807e-03 lketa = 4.336838064e-09 wketa = -1.734723476e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.735579725e-01 lpclm = 6.133304993e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.126186139e-03 lpdiblc2 = 5.474800142e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.083836002e+08 lpscbe1 = -3.362482644e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.149808009e-01 lkt1 = -1.435540156e-8
+ kt2 = -4.271211613e-02 lkt2 = 2.207348643e-9
+ at = 1.650342857e+05 lat = -1.004071626e-1
+ ute = -1.941356718e+00 lute = 7.153506284e-7
+ ua1 = 2.480362285e-11 lua1 = 1.050145812e-15
+ ub1 = -2.933984465e-19 lub1 = -2.299767186e-25
+ uc1 = 9.339214374e-12 luc1 = 7.143995830e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.40 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.878870156e-01 lvth0 = 9.076684872e-8
+ k1 = 6.324218602e-01 lk1 = -1.272284831e-7
+ k2 = -5.813040379e-02 lk2 = 3.648293062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.772314921e-02 lvoff = -6.676314387e-8
+ nfactor = 3.156179117e+00 lnfactor = -7.811282609e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 3.293471619e-02 lu0 = -8.362087220e-9
+ ua = -1.005266535e-10 lua = -1.395160132e-15
+ ub = 6.003665738e-19 lub = 1.526414650e-24
+ uc = 5.322989950e-11 luc = 2.187755377e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.446262019e+04 lvsat = -8.973374201e-3
+ a0 = 2.192553109e+00 la0 = -1.257079281e-6
+ ags = -5.161411334e-03 lags = 1.265050645e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.237329338e-24 lb0 = -4.283033172e-30
+ b1 = 0.0
+ keta = 5.265098834e-02 lketa = -1.050873655e-07 wketa = 2.428612866e-23 pketa = 4.336808690e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.147456642e-01 lpclm = 7.828278159e-7
+ pdiblc1 = 1.569430821e-01 lpdiblc1 = 4.686275877e-7
+ pdiblc2 = 6.434736582e-03 lpdiblc2 = -3.188772769e-9
+ pdiblcb = -5.007590911e-02 lpdiblcb = 5.042228697e-8
+ drout = 8.632358000e-01 ldrout = -6.097423013e-7
+ pscbe1 = 1.167628731e+09 lpscbe1 = -7.559899069e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 8.893632000e-10 lalpha0 = 5.853526093e-14
+ alpha1 = 6.266162940e-01 lalpha1 = 4.491768287e-7
+ beta0 = 1.318378417e+01 lbeta0 = 1.359725332e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.900144956e-01 lkt1 = 1.365213013e-7
+ kt2 = -4.745972127e-02 lkt2 = 1.175376658e-8
+ at = 1.651035834e+05 lat = -1.005465055e-1
+ ute = -2.002144911e+00 lute = 8.375826746e-7
+ ua1 = -5.518470310e-10 lua1 = 2.209666873e-15
+ ub1 = 6.447807678e-19 lub1 = -2.116454348e-24
+ uc1 = 1.055762826e-10 luc1 = -1.220721912e-16 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.41 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.717665141e-01 lvth0 = 5.982625921e-9
+ k1 = 4.343907494e-01 lk1 = 7.293859126e-8
+ k2 = -1.228327853e-03 lk2 = -2.103289110e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.886214874e-01 ldsub = 7.214840124e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.279980756e-01 lvoff = -5.838092139e-9
+ nfactor = 1.910881874e+00 lnfactor = 4.776007576e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -4.093947403e-22 peta0 = 7.285838599e-29
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.651219250e-02 lu0 = -1.870290187e-9
+ ua = -1.362756681e-09 lua = -1.193156915e-16
+ ub = 2.121020299e-18 lub = -1.064084691e-26
+ uc = 7.392291647e-11 luc = 9.613419190e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.218575020e+03 lvsat = 6.708225324e-2
+ a0 = 3.858874119e-01 la0 = 5.690731124e-7
+ ags = 1.309717248e+00 lags = -6.401029598e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.740171369e-02 lketa = 1.626022499e-08 wketa = -1.110223025e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.388993454e+00 lpclm = -5.051640103e-7
+ pdiblc1 = 7.437409158e-01 lpdiblc1 = -1.244994474e-7
+ pdiblc2 = 5.513544990e-03 lpdiblc2 = -2.257645204e-9
+ pdiblcb = 2.515181822e-02 lpdiblcb = -2.561684662e-08 wpdiblcb = -1.084202172e-23 ppdiblcb = 8.673617380e-30
+ drout = -4.959632800e-01 ldrout = 7.641170999e-7
+ pscbe1 = 3.120813611e+07 lpscbe1 = 3.926881210e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.191024846e-06 lalpha0 = 3.284877457e-12 walpha0 = 1.270549421e-27
+ alpha1 = 1.296767412e+00 lalpha1 = -2.282025393e-7
+ beta0 = 1.096473529e+01 lbeta0 = 3.602708867e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.301935511e-01 lkt1 = -2.502347200e-8
+ kt2 = -3.471653443e-02 lkt2 = -1.126868269e-9
+ at = 8.507713903e+04 lat = -1.965689587e-2
+ ute = -1.092230678e+00 lute = -8.214589253e-8
+ ua1 = 2.239590862e-09 lua1 = -6.118794686e-16
+ ub1 = -2.337858579e-18 lub1 = 8.983557464e-25 wub1 = -3.081487911e-39
+ uc1 = -8.386929930e-11 luc1 = 6.941675076e-17 wuc1 = 5.169878828e-32 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.42 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.215768093e-01 lvth0 = -1.945977550e-8
+ k1 = 3.667703539e-01 lk1 = 1.074781426e-7
+ k2 = 1.756159980e-02 lk2 = -3.063052309e-08 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 7.575464332e-02 ldsub = 1.297992051e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.335627272e-01 lvoff = -2.995746010e-9
+ nfactor = 2.533949421e+00 lnfactor = 1.593465777e-7
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 3.104053217e-02 lu0 = -4.183302695e-9
+ ua = -1.085244136e-09 lua = -2.610652142e-16
+ ub = 1.941064728e-18 lub = 8.127793964e-26
+ uc = 7.725809959e-11 luc = -7.422229282e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.854301274e+04 lvsat = 2.656444100e-2
+ a0 = 1.5
+ ags = 2.399526108e+00 lags = -6.206694043e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.102885254e-02 lketa = -2.318523268e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.820641385e-01 lpclm = -4.191721304e-8
+ pdiblc1 = 8.594644286e-01 lpdiblc1 = -1.836093976e-7
+ pdiblc2 = -4.584242403e-04 lpdiblc2 = 7.927530709e-10
+ pdiblcb = 1.836288000e-01 lpdiblcb = -1.065646702e-07 wpdiblcb = 1.110223025e-22 ppdiblcb = -5.551115123e-29
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.177411360e-06 lalpha0 = 3.196940107e-14
+ alpha1 = 0.85
+ beta0 = 1.686115330e+01 lbeta0 = 5.909010965e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.134635824e-01 lkt1 = 1.750969425e-8
+ kt2 = -5.758888667e-02 lkt2 = 1.055600904e-8
+ at = 7.152581445e+04 lat = -1.273506899e-2
+ ute = -2.267519941e+00 lute = 5.181754085e-7
+ ua1 = -3.630814747e-10 lua1 = 7.175291234e-16
+ ub1 = 3.233485706e-19 lub1 = -4.609516086e-25 pub1 = -3.851859889e-46
+ uc1 = 5.335421127e-11 luc1 = -6.750973096e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.43 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 7.248237971e-01 lvth0 = -4.638514448e-08 wvth0 = -2.394712385e-07 pvth0 = 6.245074640e-14
+ k1 = 4.295684749e-01 lk1 = 9.110127180e-8
+ k2 = 1.435086712e-01 lk2 = -6.347575604e-08 wk2 = -1.533740585e-07 pk2 = 3.999780722e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.865102111e-01 ldsub = -8.163449643e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.452502183e-02 lcdscd = -2.379677943e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 2.523976002e-02 lvoff = -4.440921144e-8
+ nfactor = -1.535733464e+00 lnfactor = 1.220662899e-06 wnfactor = 1.453221104e-05 pnfactor = -3.789797188e-12
+ eta0 = 1.823610115e+00 leta0 = -3.477868474e-7
+ etab = 1.175887311e-01 letab = -3.082848608e-08 petab = -4.336808690e-30
+ u0 = -5.000498844e-02 lu0 = 1.695223444e-08 wu0 = 4.063791962e-08 pu0 = -1.059780050e-14
+ ua = -4.324870790e-09 lua = 5.837840623e-16 wua = -6.692985545e-16 pua = 1.745436928e-22
+ ub = 1.603646406e-18 lub = 1.692719142e-25 wub = 3.889697840e-24 pub = -1.014378741e-30
+ uc = -1.902958301e-10 luc = 6.903209619e-17 wuc = 4.594129313e-16 puc = -1.198084607e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.974749511e+05 lvsat = -1.843483487e-03 wvsat = -9.136585120e-02 pvsat = 2.382693487e-8
+ a0 = 1.5
+ ags = -3.334129838e+00 lags = 8.745877952e-07 wags = 1.554312234e-21 pags = -8.326672685e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.455082892e-01 lketa = 1.057719111e-07 wketa = 4.665307035e-07 pketa = -1.216646760e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.154275872e-01 lpclm = -7.669653339e-08 wpclm = 3.105476395e-07 ppclm = -8.098647672e-14
+ pdiblc1 = -3.939770822e-01 lpdiblc1 = 1.432706002e-7
+ pdiblc2 = -1.329380080e-02 lpdiblc2 = 4.140039583e-09 ppdiblc2 = 3.469446952e-30
+ pdiblcb = -5.567066175e-01 lpdiblcb = 8.650444195e-8
+ drout = 2.353690284e+00 ldrout = -3.530234743e-7
+ pscbe1 = 8.233852396e+08 lpscbe1 = -6.098543103e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.221243171e-05 lalpha0 = -2.324237417e-12
+ alpha1 = 0.85
+ beta0 = 3.294674335e+01 lbeta0 = -3.603995590e-06 wbeta0 = 1.013206002e-06 pbeta0 = -2.642299403e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 6.837569132e-03 lkt1 = -6.602036187e-08 wkt1 = -5.066030008e-07 pkt1 = 1.321149702e-13
+ kt2 = 1.496186997e-02 lkt2 = -8.364212580e-9
+ at = -8.095366830e+04 lat = 2.702944539e-2
+ ute = 2.549898990e+00 lute = -7.381400046e-7
+ ua1 = 8.962747083e-09 lua1 = -1.714516403e-15
+ ub1 = -7.309374636e-18 lub1 = 1.529555746e-24
+ uc1 = -2.120305980e-10 luc1 = 6.853354557e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.44 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.816972340e-01 wvth0 = 8.786277135e-8
+ k1 = 0.90707349
+ k2 = -1.891979008e-01 wk2 = 5.627343775e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = 4.862340286e+00 wnfactor = -5.331915197e-6
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 3.884972020e-02 wu0 = -1.491018404e-8
+ ua = -1.264981373e-09 wua = 2.455678028e-16
+ ub = 2.490880869e-18 wub = -1.427142709e-24
+ uc = 1.715341584e-10 wuc = -1.685600893e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.878123790e+05 wvsat = 3.352242609e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.088925112e-01 wketa = -1.711716229e-7
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.134246447e-01 wpclm = -1.139409326e-7
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.405649150e+01 wbeta0 = -3.717485566e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.392064900e-01 wkt1 = 1.858742783e-7
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.45 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.171504489e-01 lvth0 = -1.631718124e-07 wvth0 = 4.720315981e-09 pvth0 = 3.296096131e-13
+ k1 = 4.555796457e-01 lk1 = 6.197035863e-06 wk1 = 1.329169773e-07 pk1 = -9.384885502e-12
+ k2 = 6.474164105e-03 lk2 = -2.592850776e-06 wk2 = -5.341824451e-08 pk2 = 3.948676993e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.018345153e-01 lvoff = 2.328226721e-07 wvoff = -2.874894333e-09 pvoff = -4.315619939e-13
+ nfactor = 3.068193461e+00 lnfactor = -5.376638958e-05 wnfactor = -9.389192773e-07 pnfactor = 8.357530486e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.091953141e-02 lu0 = 1.864391935e-07 wu0 = 1.118635428e-09 pu0 = -3.112530291e-13
+ ua = -7.558861509e-10 lua = -1.482132562e-15 wua = 4.467832666e-17 pua = 3.012020984e-21
+ ub = 1.549535476e-18 lub = 1.380658775e-23 wub = -2.760243305e-26 pub = -2.415799785e-29
+ uc = -7.319592212e-11 luc = 5.364165217e-15 wuc = 1.790877147e-16 puc = -7.480901143e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.090524119e+00 la0 = 1.129571087e-05 wa0 = 4.310059281e-07 pa0 = -1.521223700e-11
+ ags = 3.090914179e-01 lags = 4.137844151e-06 wags = 1.099036507e-07 pags = -6.054113547e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.198190121e-24 lb0 = 3.418877166e-28 wb0 = 1.363034970e-29 pb0 = -4.545573362e-34
+ b1 = 0.0
+ keta = -5.303646030e-03 lketa = -2.334581660e-07 wketa = -1.596515128e-09 pketa = 3.877846151e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.242116906e-02 lpclm = 6.225321695e-07 wpclm = 3.583640978e-08 ppclm = -7.171147271e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 6.355388330e-03 lpdiblc2 = -1.156498144e-07 wpdiblc2 = -4.682491401e-09 ppdiblc2 = 1.530420327e-13
+ pdiblcb = 9.324003944e+00 lpdiblcb = -2.529245211e-04 wpdiblcb = -1.371827341e-05 ppdiblcb = 2.997970971e-10
+ drout = 0.56
+ pscbe1 = 3.084204719e+08 lpscbe1 = 1.146351867e+04 wpscbe1 = 5.680178049e+02 ppscbe1 = -1.412739309e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.376827215e-01 lkt1 = -8.824353779e-07 wkt1 = 1.771038384e-08 pkt1 = 1.704077709e-12
+ kt2 = -4.786010220e-02 lkt2 = -9.849535387e-07 wkt2 = 1.946113545e-09 pkt2 = 1.723185705e-12
+ at = 140000.0
+ ute = -1.882501289e+00 lute = -2.573942053e-05 wute = -3.860869844e-08 pute = 4.413345560e-11
+ ua1 = 6.966609528e-10 lua1 = -6.345000468e-14 wua1 = -7.160395961e-16 pua1 = 1.025617504e-19
+ ub1 = -1.119883260e-18 lub1 = 4.227123315e-23 wub1 = 9.492126458e-25 pub1 = -6.358906180e-29
+ uc1 = -3.282482510e-12 luc1 = 2.541245255e-15 wuc1 = 3.265619405e-17 puc1 = -4.067790957e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.46 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.089962558e-01 wvth0 = 2.119191350e-8
+ k1 = 7.652644259e-01 wk1 = -3.360743707e-7
+ k2 = -1.230984961e-01 wk2 = 1.439091864e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.019965643e-02 wvoff = -2.444136323e-8
+ nfactor = 3.813230110e-01 wnfactor = 3.237593572e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.023646647e-02 wu0 = -1.443562762e-8
+ ua = -8.299528348e-10 wua = 1.951982005e-16
+ ub = 2.239492770e-18 wub = -1.234851256e-24
+ uc = 1.948677720e-10 wuc = -1.947557287e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.655005238e+00 wa0 = -3.291959449e-7
+ ags = 5.158721086e-01 wags = -1.926388654e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.886981675e-24 wb0 = -9.085266575e-30
+ b1 = 0.0
+ keta = -1.697026253e-02 wketa = 1.778226465e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 5.760144238e-04 wpdiblc2 = 2.965485678e-9
+ pdiblcb = -3.315405677e+00 wpdiblcb = 1.263501771e-6
+ drout = 0.56
+ pscbe1 = 8.812874582e+08 wpscbe1 = -1.379711096e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.817807084e-01 wkt1 = 1.028683436e-7
+ kt2 = -9.708123418e-02 wkt2 = 8.805895814e-8
+ at = 140000.0
+ ute = -3.168778627e+00 wute = 2.166874665e-6
+ ua1 = -2.474129274e-09 wua1 = 4.409283838e-15
+ ub1 = 9.925391686e-19 wub1 = -2.228526689e-24
+ uc1 = 1.237112925e-10 wuc1 = -1.706237249e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.47 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910522174e-01 lvth0 = 1.437458519e-07 wvth0 = 2.997572762e-08 pvth0 = -7.036525518e-14
+ k1 = 7.994523375e-01 lk1 = -2.738720441e-07 wk1 = -3.947886715e-07 pk1 = 4.703476985e-13
+ k2 = -1.351107206e-01 lk2 = 9.622735951e-08 wk2 = 1.684724982e-07 pk2 = -1.967714338e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -8.299661719e-02 lvoff = -5.770200590e-08 wvoff = -3.898426245e-08 pvoff = 1.165000535e-13
+ nfactor = 1.858059204e-01 lnfactor = 1.566245571e-06 wnfactor = 3.782761542e-06 pnfactor = -4.367223944e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.891653727e-02 lu0 = 1.057367036e-08 wu0 = -1.244101576e-08 pu0 = -1.597840875e-14
+ ua = -9.813544586e-10 lua = 1.212846008e-15 wua = 4.137751516e-16 pua = -1.750973179e-21
+ ub = 2.304602062e-18 lub = -5.215766049e-25 wub = -1.321137456e-24 pub = 6.912202832e-31
+ uc = 2.324585165e-10 luc = -3.011314097e-16 wuc = -2.375702840e-16 puc = 3.429782407e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.513699368e+00 la0 = 1.131971079e-06 wa0 = -1.427725248e-08 pa0 = -2.522746252e-12
+ ags = 3.813023510e-01 lags = 1.078009531e-06 wags = -2.665599029e-08 pags = -1.329653292e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.579523060e-23 lb0 = -6.335128974e-29 wb0 = -1.819503157e-29 pb0 = 7.297637790e-35
+ b1 = 0.0
+ keta = -4.569511354e-03 lketa = -9.933976387e-08 wketa = -9.546900219e-09 pketa = 2.189280913e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.010244142e-01 lpclm = 2.279512528e-06 wpclm = -1.915501765e-07 ppclm = 1.534467472e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.750100865e-03 lpdiblc2 = 2.664479779e-08 wpdiblc2 = 6.572556201e-09 ppdiblc2 = -2.889547005e-14
+ pdiblcb = -6.614683933e+00 lpdiblcb = 2.642981206e-05 wpdiblcb = 2.530410575e-06 ppdiblcb = -1.014893531e-11
+ drout = 0.56
+ pscbe1 = 8.121675033e+08 lpscbe1 = 5.537051663e+02 wpscbe1 = -3.953947846e+01 ppscbe1 = -7.885147326e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.768321321e-01 lkt1 = -3.964198524e-08 wkt1 = 9.858861725e-08 pkt1 = 3.428397196e-14
+ kt2 = -9.312253560e-02 lkt2 = -3.171228714e-08 wkt2 = 8.357010014e-08 pkt2 = 3.595928076e-14
+ at = 140000.0
+ ute = -2.715161340e+00 lute = -3.633831010e-06 wute = 1.410789675e-06 pute = 6.056835047e-12
+ ua1 = -2.027849365e-09 lua1 = -3.575052845e-15 wua1 = 3.777501339e-15 pua1 = 5.061074396e-21
+ ub1 = 6.961711965e-19 lub1 = 2.374140402e-24 wub1 = -1.879958151e-24 pub1 = -2.792307964e-30
+ uc1 = 9.557869579e-11 luc1 = 2.253642120e-16 wuc1 = -1.452897767e-16 puc1 = -2.029448378e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.48 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.078368527e-01 lvth0 = -3.246523284e-07 wvth0 = -1.120050086e-07 pvth0 = 4.990890939e-13
+ k1 = 8.120910460e-01 lk1 = -3.245631992e-07 wk1 = -4.276800911e-07 pk1 = 6.022681437e-13
+ k2 = -1.644818103e-01 lk2 = 2.140285150e-07 wk2 = 2.109338787e-07 pk2 = -3.670749443e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.625454835e-01 lvoff = 2.613514734e-07 wvoff = 8.810008177e-08 pvoff = -3.932080551e-13
+ nfactor = -2.962307874e+00 lnfactor = 1.419265630e-05 wnfactor = 7.501482573e-06 pnfactor = -1.928221819e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.471392842e-02 lu0 = -1.267842493e-08 wu0 = -1.771484690e-08 pu0 = 5.173799349e-15
+ ua = -1.553357880e-09 lua = 3.507029322e-15 wua = 1.511181270e-15 pua = -6.152434275e-21
+ ub = 3.913268596e-18 lub = -6.973593817e-24 wub = -3.748765726e-24 pub = 1.042791776e-29
+ uc = 2.235302459e-10 luc = -2.653220272e-16 wuc = -2.615174968e-16 puc = 4.390253863e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 3.535560920e-01 la0 = 5.785057490e-06 wa0 = 1.338507215e-06 pa0 = -7.948475256e-12
+ ags = 4.463057386e-01 lags = 8.172948537e-07 wags = -3.567002700e-07 pags = -5.916316050e-15
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.929516167e-24 lb0 = 3.180359243e-29 wb0 = 9.134263418e-30 pb0 = -3.663557584e-35
+ b1 = 0.0
+ keta = -8.468260840e-02 lketa = 2.219767242e-07 wketa = 1.303367018e-07 pketa = -3.421151014e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.760744296e-01 lpclm = -3.510743488e-08 wpclm = 1.532375006e-07 ppclm = 1.515978842e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 4.167704910e-03 lpdiblc2 = -1.101040765e-09 wpdiblc2 = -3.209128685e-09 ppdiblc2 = 1.033677475e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.132630470e+09 lpscbe1 = -7.316032133e+02 wpscbe1 = -5.096940303e+02 ppscbe1 = 1.097174562e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.677224275e-01 lkt1 = -7.617906097e-08 wkt1 = 8.290625060e-08 pkt1 = 9.718258858e-14
+ kt2 = -9.481774513e-02 lkt2 = -2.491316450e-08 wkt2 = 8.190650560e-08 pkt2 = 4.263160247e-14
+ at = 1.542800880e+05 lat = -5.727437697e-02 wat = 1.690486752e-02 pat = -6.780180599e-8
+ ute = -2.460414528e+00 lute = -4.655565958e-06 wute = 8.159235804e-07 pute = 8.442715652e-12
+ ua1 = 2.043774588e-09 lua1 = -1.990546520e-14 wua1 = -3.173685068e-15 pua1 = 3.294079552e-20
+ ub1 = -3.427478360e-18 lub1 = 1.891321631e-23 wub1 = 4.926560507e-24 pub1 = -3.009179771e-29
+ uc1 = 5.219392052e-11 luc1 = 3.993712613e-16 wuc1 = -6.736468393e-17 puc1 = -5.154857089e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.49 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 3.607891851e-01 lvth0 = 1.721076630e-07 wvth0 = 1.997891469e-07 pvth0 = -1.278622288e-13
+ k1 = 7.207257604e-01 lk1 = -1.408471619e-07 wk1 = -1.388077264e-07 pk1 = 2.140763709e-14
+ k2 = -7.661043593e-02 lk2 = 3.733798554e-08 wk2 = 2.904935389e-08 pk2 = -1.344088184e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 2.102585095e-02 lvoff = -1.077711959e-07 wvoff = -1.395073933e-07 pvoff = 6.446186923e-14
+ nfactor = 4.244063249e+00 lnfactor = -2.978138602e-07 wnfactor = -1.710079880e-06 pnfactor = -7.597373725e-13
+ eta0 = 1.583044666e-01 leta0 = -1.574535251e-07 weta0 = -2.178916211e-13 peta0 = 4.381334211e-19
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 4.680736892e-02 lu0 = -1.688788579e-08 wu0 = -2.180686675e-08 pu0 = 1.340197559e-14
+ ua = 2.141002321e-09 lua = -3.921538449e-15 wua = -3.523531124e-15 pua = 3.971294921e-21
+ ub = -1.868587428e-18 lub = 4.652481330e-24 wub = 3.881027802e-24 pub = -4.913964248e-30
+ uc = 9.535499624e-11 luc = -7.589029566e-18 wuc = -6.621778757e-17 puc = 4.631946528e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.244250068e+05 lvsat = -8.932918177e-02 wvsat = -6.281815435e-02 pvsat = 1.263138653e-7
+ a0 = 4.283641088e+00 la0 = -2.117502399e-06 wa0 = -3.287048110e-06 pa0 = 1.352526634e-12
+ ags = -1.023502674e+00 lags = 3.772765031e-06 wags = 1.600763217e-06 pags = -3.941956491e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.585903233e-23 lb0 = -1.603008786e-29 wb0 = -1.826852684e-29 pb0 = 1.846557117e-35
+ b1 = 0.0
+ keta = 2.722724700e-01 lketa = -4.957835501e-07 wketa = -3.452300349e-07 pketa = 6.141478349e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.346917266e-01 lpclm = 2.198405601e-06 wpclm = 1.335257817e-06 ppclm = -2.225192019e-12
+ pdiblc1 = -6.244660677e-01 lpdiblc1 = 2.039874166e-06 wpdiblc1 = 1.228322048e-06 ppdiblc1 = -2.469892777e-12
+ pdiblc2 = 1.096863474e-02 lpdiblc2 = -1.477625526e-08 wpdiblc2 = -7.126979603e-09 ppdiblc2 = 1.821473452e-14
+ pdiblcb = -1.864189408e-01 lpdiblcb = 3.245789463e-07 wpdiblcb = 2.143219745e-07 ppdiblcb = -4.309556259e-13
+ drout = 1.243869036e+00 ldrout = -1.375114283e-06 wdrout = -5.983295634e-07 pdrout = 1.203112709e-12
+ pscbe1 = 2.175922303e+09 lpscbe1 = -2.829439825e+03 wpscbe1 = -1.584968930e+03 ppscbe1 = 3.259322276e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.227897527e-08 lalpha0 = 2.257689916e-13 walpha0 = 1.307349726e-13 palpha0 = -2.628800527e-19
+ alpha1 = -4.102156589e-01 lalpha1 = 2.534024004e-06 walpha1 = 1.629829325e-06 palpha1 = -3.277237990e-12
+ beta0 = 1.132913022e+01 lbeta0 = 5.089037525e-06 wbeta0 = 2.915389890e-06 pbeta0 = -5.862225174e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.625754292e-01 lkt1 = 3.156286268e-07 wkt1 = 2.712540534e-07 pkt1 = -2.815445364e-13
+ kt2 = -1.804497844e-01 lkt2 = 1.472745412e-07 wkt2 = 2.090513359e-07 pkt2 = -2.130294423e-13
+ at = 2.422931815e+05 lat = -2.342498731e-01 wat = -1.213367992e-01 pat = 2.101726021e-7
+ ute = -8.065528057e+00 lute = 6.615117856e-06 wute = 9.531225997e-06 pute = -9.081892433e-12
+ ua1 = -1.852321893e-08 lua1 = 2.145035744e-14 wua1 = 2.824977458e-14 pua1 = -3.024505721e-20
+ ub1 = 1.537495432e-17 lub1 = -1.889445208e-23 wub1 = -2.315483117e-23 pub1 = 2.637387153e-29
+ uc1 = 6.118300250e-10 luc1 = -7.259371827e-16 wuc1 = -7.957964577e-16 puc1 = 9.492347038e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.50 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.006127632e-01 lvth0 = 3.077594773e-08 wvth0 = 1.118488580e-07 pvth0 = -3.897341593e-14
+ k1 = 5.472829464e-01 lk1 = 3.446640629e-08 wk1 = -1.774588569e-07 pk1 = 6.047565865e-14
+ k2 = -2.083649143e-02 lk2 = -1.903753673e-08 wk2 = 3.082269978e-08 pk2 = -3.136561385e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.423481142e-01 ldsub = 1.189208791e-07 wdsub = 7.273859612e-08 pdsub = -7.352315462e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -4.744689245e-02 lvoff = -3.855990548e-08 wvoff = -1.266209824e-07 pvoff = 5.143646549e-14
+ nfactor = 5.440351800e+00 lnfactor = -1.507005579e-06 wnfactor = -5.548086719e-06 pnfactor = 3.119666208e-12
+ eta0 = -4.954534531e-01 leta0 = 5.033558275e-07 weta0 = 4.357832419e-13 peta0 = -2.225919791e-19
+ etab = -1.690560735e-01 letab = 8.559444360e-08 wetab = -1.376354510e-09 petab = 1.391199869e-15
+ u0 = 3.385321651e-02 lu0 = -3.794009886e-09 wu0 = -1.153959056e-08 pu0 = 3.023956554e-15
+ ua = -1.573012728e-09 lua = -1.674640342e-16 wua = 3.305082081e-16 pua = 7.568592061e-23
+ ub = 2.487104708e-18 lub = 2.498086988e-25 wub = -5.754597958e-25 pub = -4.094089753e-31
+ uc = 1.050098941e-10 luc = -1.734806517e-17 wuc = -4.886661494e-17 puc = 2.878114290e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.943727398e+04 lvsat = 8.640837759e-02 wvsat = 9.220300603e-02 pvsat = -3.037935331e-8
+ a0 = 2.892326084e+00 la0 = -7.111806710e-07 wa0 = -3.939951154e-06 pa0 = 2.012471890e-12
+ ags = 4.016569868e+00 lags = -1.321669733e-06 wags = -4.254988253e-06 pags = 1.976955114e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.938196835e-01 lketa = 1.774930733e-07 wketa = 5.131068521e-07 pketa = -2.534470738e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.783136245e+00 lpclm = -1.357365663e-06 wpclm = -2.191497666e-06 ppclm = 1.339603049e-12
+ pdiblc1 = 1.303826661e+00 lpdiblc1 = 9.078287259e-08 wpdiblc1 = -8.804167052e-07 ppdiblc1 = -3.384091679e-13
+ pdiblc2 = -7.060664760e-03 lpdiblc2 = 3.447508269e-09 wpdiblc2 = 1.976580268e-08 ppdiblc2 = -8.968113309e-15
+ pdiblcb = 2.978378816e-01 lpdiblcb = -1.649010702e-07 wpdiblcb = -4.286439490e-07 ppdiblcb = 2.189453282e-13
+ drout = -1.257229751e+00 ldrout = 1.152961356e-06 wdrout = 1.196659127e-06 pdrout = -6.112367287e-13
+ pscbe1 = -2.077353648e+09 lpscbe1 = 1.469711960e+03 wpscbe1 = 3.314515743e+03 ppscbe1 = -1.693008238e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.201866089e-05 lalpha0 = 1.229089672e-11 walpha0 = 1.387644358e-11 palpha0 = -1.415684987e-17
+ alpha1 = 3.370431318e+00 lalpha1 = -1.287401031e-06 walpha1 = -3.259658651e-06 palpha1 = 1.664988004e-12
+ beta0 = 3.023906564e+00 lbeta0 = 1.348384132e-05 wbeta0 = 1.248244278e-05 pbeta0 = -1.553246830e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.972282506e-01 lkt1 = -5.365918644e-08 wkt1 = -5.181921065e-08 pkt1 = 4.501339586e-14
+ kt2 = -3.092003953e-02 lkt2 = -3.868031485e-09 wkt2 = -5.967831825e-09 pkt2 = 4.308922176e-15
+ at = -1.637544366e+04 lat = 2.720875177e-02 wat = 1.594765612e-01 pat = -7.366961124e-8
+ ute = -1.718773352e+00 lute = 1.999070543e-07 wute = 9.848824781e-07 pute = -4.433680528e-13
+ ua1 = 4.536080362e-09 lua1 = -1.857659456e-15 wua1 = -3.609925333e-15 pua1 = 1.958281428e-21
+ ub1 = -6.397761641e-18 lub1 = 3.113104392e-24 wub1 = 6.381891540e-24 pub1 = -3.481434268e-30
+ uc1 = -3.041207366e-10 luc1 = 1.998930238e-16 wuc1 = 3.462202823e-16 puc1 = -2.050998288e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.51 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.086461845e-01 lvth0 = -2.440601139e-08 wvth0 = 2.032606287e-08 pvth0 = 7.775146479e-15
+ k1 = 8.102388335e-01 lk1 = -9.984777950e-08 wk1 = -6.971022941e-07 pk1 = 3.259022514e-13
+ k2 = -1.499352824e-01 lk2 = 4.690431832e-08 wk2 = 2.632937091e-07 pk2 = -1.218794983e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.602808753e-01 ldsub = 2.734995301e-07 wdsub = 3.710317849e-07 pdsub = -2.258871393e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -4.178715321e-03 lcdscd = 4.892673684e-09 wcdscd = 1.505708913e-08 pcdscd = -7.690950329e-15
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.955161298e-01 lvoff = 3.707178801e-08 wvoff = 9.738653616e-08 pvoff = -6.298343888e-14
+ nfactor = -2.910502403e+00 lnfactor = 2.758493836e-06 wnfactor = 8.558308045e-06 pnfactor = -4.085682748e-12
+ eta0 = -9.099168273e-01 leta0 = 7.150579165e-07 weta0 = 2.200574058e-06 peta0 = -1.124022421e-12
+ etab = -1.264674471e-01 letab = 6.384076948e-08 wetab = 1.978157696e-07 petab = -1.003533484e-13
+ u0 = 4.874596896e-02 lu0 = -1.140101934e-08 wu0 = -2.783174266e-08 pu0 = 1.134575976e-14
+ ua = 1.098853166e-09 lua = -1.532215726e-15 wua = -3.433252440e-15 pua = 1.998162167e-21
+ ub = 1.624399029e-19 lub = 1.437214936e-24 wub = 2.795877278e-24 pub = -2.131440754e-30
+ uc = 1.194575444e-10 luc = -2.472772268e-17 wuc = -6.633465772e-17 puc = 3.770357460e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.239741596e+04 lvsat = 1.906906366e-02 wvsat = 9.660460239e-03 pvsat = 1.178222349e-8
+ a0 = 1.5
+ ags = 6.419781951e+00 lags = -2.549196820e-06 wags = -6.319568808e-06 pags = 3.031513958e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.766946049e-01 lketa = 6.658862296e-08 wketa = 2.289766575e-07 pketa = -1.083173482e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.150865120e-01 lpclm = 2.251631461e-07 wpclm = 1.253066616e-06 ppclm = -4.198321631e-13
+ pdiblc1 = 3.441624505e+00 lpdiblc1 = -1.001174337e-06 wpdiblc1 = -4.058980054e-06 ppdiblc1 = 1.285156491e-12
+ pdiblc2 = 1.333581783e-02 lpdiblc2 = -6.970729485e-09 wpdiblc2 = -2.168361052e-08 ppdiblc2 = 1.220366666e-14
+ pdiblcb = 5.318277763e-01 lpdiblcb = -2.844198325e-07 wpdiblcb = -5.473451131e-07 ppdiblcb = 2.795762210e-13
+ drout = -4.209953797e-01 ldrout = 7.258245460e-07 wdrout = 2.233708109e-06 pdrout = -1.140946830e-12
+ pscbe1 = 7.754520529e+08 lpscbe1 = 1.253874771e+01 wpscbe1 = 3.858770358e+01 ppscbe1 = -1.971005876e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.178576889e-05 lalpha0 = 1.319272505e-13 walpha0 = -1.353175267e-11 palpha0 = -1.571269422e-19
+ alpha1 = 0.85
+ beta0 = 2.640847418e+01 lbeta0 = 1.539331569e-06 wbeta0 = -1.500773919e-05 pbeta0 = -1.490868209e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.453160813e-01 lkt1 = 2.198200426e-08 wkt1 = 5.006996227e-08 pkt1 = -7.030167216e-15
+ kt2 = -9.446450759e-02 lkt2 = 2.858959318e-08 wkt2 = 5.796596854e-08 pkt2 = -2.834756798e-14
+ at = 6.895266352e+04 lat = -1.637565078e-02 wat = 4.044818287e-03 pat = 5.722747009e-9
+ ute = -5.390597267e+00 lute = 2.075423305e-06 wute = 4.909265188e-06 pute = -2.447887800e-12
+ ua1 = -7.555439804e-09 lua1 = 4.318519763e-15 wua1 = 1.130589821e-14 pua1 = -5.660512418e-21
+ ub1 = 7.044167282e-18 lub1 = -3.752844715e-24 wub1 = -1.056467000e-23 pub1 = 5.174632115e-30
+ uc1 = 4.011161556e-10 luc1 = -1.603321074e-16 wuc1 = -5.466581287e-16 puc1 = 2.509699632e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.52 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.009440125e-01 lvth0 = 3.681207239e-09 wvth0 = 1.124525592e-07 pvth0 = -1.625015399e-14
+ k1 = -8.800822560e-01 lk1 = 3.409642962e-07 wk1 = 2.058681893e-06 pk1 = -3.927676836e-13
+ k2 = 5.270626092e-01 lk2 = -1.296472538e-07 wk2 = -7.562947674e-07 pk2 = 1.440149021e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.060018301e+00 ldsub = -3.055234108e-07 wdsub = -1.844674918e-06 pdsub = 3.519381490e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.873471940e-02 lcdscd = -8.906409304e-09 wcdscd = -5.377531833e-08 pcdscd = 1.025957788e-14
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 3.668248164e-01 lvoff = -1.095788580e-07 wvoff = -5.369484809e-07 pvoff = 1.024422529e-13
+ nfactor = 2.625586680e+01 lnfactor = -4.847686923e-06 wnfactor = -2.915429475e-05 pnfactor = 5.749236084e-12
+ eta0 = 6.823313069e+00 leta0 = -1.301660175e-06 weta0 = -7.859193065e-06 peta0 = 1.499424008e-12
+ etab = 5.607718891e-01 letab = -1.153816281e-07 wetab = -6.966537879e-07 petab = 1.329117896e-13
+ u0 = -6.200883872e-02 lu0 = 1.748228394e-08 wu0 = 5.950715600e-08 pu0 = -1.143100227e-14
+ ua = -1.466912303e-08 lua = 2.579851715e-15 wua = 1.559116256e-14 pua = -2.963138924e-21
+ ub = 1.883521419e-17 lub = -3.432383179e-24 wub = -2.319715496e-23 pub = 4.647178152e-30
+ uc = 4.150765126e-11 luc = -4.399481842e-18 wuc = 9.503362116e-17 puc = -4.379013379e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.049693872e+05 lvsat = -1.289599042e-02 wvsat = -1.031465950e-01 pvsat = 4.120072420e-8
+ a0 = 1.5
+ ags = -1.590700091e+01 lags = 3.273315576e-06 wags = 1.976369838e-05 pags = -3.770636959e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.929877674e-01 lketa = -5.589796420e-08 wketa = -6.943348799e-07 pketa = 1.324693744e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.658623088e+00 lpclm = -2.895526856e-07 wpclm = -1.329284751e-06 ppclm = 2.536089204e-13
+ pdiblc1 = -2.453601965e+00 lpdiblc1 = 5.362181932e-07 wpdiblc1 = 3.237590262e-06 ppdiblc1 = -6.176868957e-13
+ pdiblc2 = -7.281004859e-02 lpdiblc2 = 1.549490643e-08 wpdiblc2 = 9.355549441e-08 ppdiblc2 = -1.784907856e-14
+ pdiblcb = -1.800274390e+00 lpdiblcb = 3.237597630e-07 wpdiblcb = 1.954803975e-06 ppdiblcb = -3.729492313e-13
+ drout = 7.428673782e+00 ldrout = -1.321259276e-06 wdrout = -7.977528961e-06 pdrout = 1.522000840e-12
+ pscbe1 = 9.110564793e+08 lpscbe1 = -2.282498823e+01 wpscbe1 = -1.378132271e+02 ppscbe1 = 2.629283434e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.571095995e-05 lalpha0 = -8.715287625e-12 walpha0 = -5.265740848e-11 palpha0 = 1.004629633e-17
+ alpha1 = 0.85
+ beta0 = 8.293324901e+01 lbeta0 = -1.320153836e-05 wbeta0 = -7.756218182e-05 pbeta0 = 1.482245466e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.702197084e-01 lkt1 = 2.847652154e-08 wkt1 = 8.610539949e-08 pkt1 = -1.642770475e-14
+ kt2 = 1.352038480e-01 lkt2 = -3.130469859e-08 wkt2 = -1.890122130e-07 pkt2 = 3.606088406e-14
+ at = -2.920533911e+05 lat = 7.776967419e-02 wat = 3.318344095e-01 pat = -7.976018933e-8
+ ute = 1.316122831e+01 lute = -2.762633080e-06 wute = -1.668028812e-05 pute = 3.182365449e-12
+ ua1 = 3.361023680e-08 lua1 = -6.416912376e-15 wua1 = -3.874417781e-14 pua1 = 7.391846708e-21
+ ub1 = -2.929791289e-17 lub1 = 5.724661006e-24 wub1 = 3.456448692e-23 pub1 = -6.594420202e-30
+ uc1 = -1.197252937e-09 luc1 = 2.565001747e-16 wuc1 = 1.548702521e-15 puc1 = -2.954707592e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.53 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.202389672e-01 wvth0 = 2.727778751e-8
+ k1 = 0.90707349
+ k2 = -1.524801971e-01 wk2 = -1.444295688e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = 8.468382376e-01 wnfactor = 9.801809689e-7
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 2.962411096e-02 wu0 = -4.081536500e-10
+ ua = -1.146895435e-09 wua = 5.994473803e-17
+ ub = 8.444644532e-19 wub = 1.160911940e-24
+ uc = 1.844787831e-11 wuc = 7.208113314e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.373753791e+05 wvsat = 1.128059602e-1
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 0.0
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.14094
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.373771914e+01 wbeta0 = 1.293399123e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 1.155743918e+05 wat = -8.622660822e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.54 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.984260027e-01 lvth0 = -3.422502814e-06 wvth0 = -2.040967952e-07 pvth0 = 4.084137293e-12
+ k1 = 5.000310512e-01 lk1 = -5.305874165e-07 wk1 = 8.171198085e-08 pk1 = -1.635120962e-12
+ k2 = -3.823891573e-02 lk2 = 8.018114364e-07 wk2 = -1.911817029e-09 pk2 = 3.825696143e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.348192401e-02 lvoff = -3.589023715e-07 wvoff = -1.249651158e-08 pvoff = 2.500650189e-13
+ nfactor = -4.099373251e+00 lnfactor = 1.459041087e-04 wnfactor = 7.317630180e-06 pnfactor = -1.464315316e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.069728418e-02 lu0 = -8.603134005e-07 wu0 = -4.470263087e-08 pu0 = 8.945347799e-13
+ ua = 7.554738052e-10 lua = -2.833474780e-14 wua = -1.696305570e-15 pua = 3.394440776e-20
+ ub = 2.407223415e-18 lub = -2.480763985e-23 wub = -1.015600616e-24 pub = 2.032296659e-29
+ uc = 1.784860171e-10 luc = -3.055387225e-15 wuc = -1.108327650e-16 puc = 2.217850741e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.820568239e+00 la0 = -9.031672940e-06 wa0 = -4.099552559e-07 pa0 = 8.203526896e-12
+ ags = 6.122520352e-01 lags = -5.275064012e-06 wags = -2.393167654e-07 pags = 4.788916579e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.134409340e-08 lb0 = -1.227543525e-12 wb0 = -7.066422420e-14 pb0 = 1.414046668e-18
+ b1 = -5.307138953e-08 lb1 = 1.062000219e-12 wb1 = 6.113463188e-14 pb1 = -1.223352036e-18
+ keta = -1.145550966e-02 lketa = 1.985500596e-07 wketa = 5.490013447e-09 pketa = -1.098594842e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.693917305e-01 lpclm = -5.720297905e-06 wpclm = -3.292921230e-07 ppclm = 6.589394206e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 8.732858526e-03 lpdiblc2 = -1.117099292e-07 wpdiblc2 = -7.421175400e-09 ppdiblc2 = 1.485035528e-13
+ pdiblcb = -1.324901929e+01 lpdiblcb = 2.207283363e-04 wpdiblcb = 1.228431438e-05 ppdiblcb = -2.458187862e-10
+ drout = 0.56
+ pscbe1 = 3.239655734e+09 lpscbe1 = -4.958956792e+04 wpscbe1 = -2.808565893e+03 ppscbe1 = 5.620161106e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.507945870e-01 lkt1 = 3.167999322e-06 wkt1 = 1.480075613e-07 pkt1 = -2.961747636e-12
+ kt2 = -9.567707948e-02 lkt2 = 1.501617896e-06 wkt2 = 5.702801982e-08 pkt2 = -1.141175501e-12
+ at = -1.010089968e+04 lat = 3.003636982e+00 wat = 1.729060296e-01 pat = -3.459985556e-6
+ ute = -4.810391969e+00 lute = 7.049183513e-05 wute = 3.334122267e-06 pute = -6.671840719e-11
+ ua1 = -3.313444255e-09 lua1 = 9.339122385e-14 wua1 = 3.903328917e-15 pua1 = -7.810867964e-20
+ ub1 = 3.230221434e-19 lub1 = -2.531528804e-23 wub1 = -7.129162608e-25 pub1 = 1.426601473e-29
+ uc1 = -5.492017226e-11 luc1 = 6.105660860e-16 wuc1 = 9.213930127e-17 puc1 = -1.843779840e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.55 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.5273931
+ k1 = 0.47351598
+ k2 = 0.0018300469
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.11141737
+ nfactor = 3.1919
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0277048
+ ua = -6.6049995e-10
+ ub = 1.16751e-18
+ uc = 2.5799e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.369228
+ ags = 0.348641
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0015333577
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0031503727
+ pdiblcb = -2.2185512
+ drout = 0.56
+ pscbe1 = 761513800.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.29248
+ kt2 = -0.020636654
+ at = 140000.0
+ ute = -1.2877
+ ua1 = 1.3536e-9
+ ub1 = -9.4206e-19
+ uc1 = -2.4408323e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.56 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.170743503e-01 lvth0 = 8.266129549e-8
+ k1 = 4.567336080e-01 lk1 = 1.344399904e-7
+ k2 = 1.114140034e-02 lk2 = -7.459125980e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.168391204e-01 lvoff = 4.343248247e-8
+ nfactor = 3.469646931e+00 lnfactor = -2.224971222e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.811640691e-02 lu0 = -3.297294898e-9
+ ua = -6.221534367e-10 lua = -3.071857119e-16
+ ub = 1.157713655e-18 lub = 7.847642182e-26
+ uc = 2.622213792e-11 luc = -3.389667350e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.501305188e+00 la0 = -1.058042092e-6
+ ags = 3.581621046e-01 lags = -7.627153156e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.285724033e-02 lketa = 9.071320047e-08 wketa = -1.734723476e-24 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.673104246e-01 lpclm = 3.611594172e-06 wpclm = 1.110223025e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 2.955579854e-03 lpdiblc2 = 1.560443807e-9
+ pdiblcb = -4.418017311e+00 lpdiblcb = 1.761945233e-5
+ drout = 0.56
+ pscbe1 = 7.778430133e+08 lpscbe1 = -1.308098334e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912466833e-01 lkt1 = -9.879836114e-9
+ kt2 = -2.057476356e-02 lkt2 = -4.957910604e-10
+ at = 140000.0
+ ute = -1.490445232e+00 lute = 1.624148668e-6
+ ua1 = 1.251425227e-09 lua1 = 8.185002439e-16
+ ub1 = -9.358332547e-19 lub1 = -4.988112379e-26
+ uc1 = -3.054834705e-11 luc1 = 4.918641870e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.57 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.106045433e-01 lvth0 = 1.086103068e-7
+ k1 = 4.408190516e-01 lk1 = 1.982698706e-7
+ k2 = 1.863132370e-02 lk2 = -1.046317395e-07 wk2 = 6.938893904e-24
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -8.606520361e-02 lvoff = -7.999511228e-8
+ nfactor = 3.549780143e+00 lnfactor = -2.546368387e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.933554941e-02 lu0 = -8.187014548e-9
+ ua = -2.414911465e-10 lua = -1.833940696e-15
+ ub = 6.589395849e-19 lub = 2.078952480e-24
+ uc = -3.494870781e-12 luc = 1.157988951e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.515523305e+00 la0 = -1.115067914e-6
+ ags = 1.366518094e-01 lags = 8.121588595e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.846356849e-02 lketa = -7.501572108e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.091009455e-01 lpclm = 9.649571892e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.381838483e-03 lpdiblc2 = 7.872383663e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.901616173e+08 lpscbe1 = 2.208614822e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957509478e-01 lkt1 = 8.185804823e-9
+ kt2 = -2.371415082e-02 lkt2 = 1.209561941e-8
+ at = 1.689553184e+05 lat = -1.161335857e-1
+ ute = -1.752105721e+00 lute = 2.673612892e-6
+ ua1 = -7.113229936e-10 lua1 = 8.690663327e-15 pua1 = 3.308722450e-36
+ ub1 = 8.493023065e-19 lub1 = -7.209677841e-24
+ uc1 = -6.285819551e-12 luc1 = -4.812538692e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.58 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.342275017e-01 lvth0 = 6.110959292e-8
+ k1 = 6.002258295e-01 lk1 = -1.222630466e-7
+ k2 = -5.139249434e-02 lk2 = 3.617117345e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.000814656e-01 lvoff = -5.181140900e-8
+ nfactor = 2.759531280e+00 lnfactor = -9.573470380e-7
+ eta0 = 1.583042774e-01 leta0 = -1.574531447e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 2.787667965e-02 lu0 = -5.253539668e-9
+ ua = -9.177990006e-10 lua = -4.740303314e-16
+ ub = 1.500559190e-18 lub = 3.866355608e-25
+ uc = 3.787088470e-11 luc = 3.262121312e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.989214000e+04 lvsat = 2.032474338e-2
+ a0 = 1.430132279e+00 la0 = -9.433648340e-7
+ ags = 3.661307571e-01 lags = 3.507258042e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.742407017e-02 lketa = 3.736236032e-08 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.244546611e-01 lpclm = 2.667012826e-7
+ pdiblc1 = 4.418486520e-01 lpdiblc1 = -1.042565435e-7
+ pdiblc2 = 4.781655300e-03 lpdiblc2 = 1.036079606e-9
+ pdiblcb = -3.645777836e-04 lpdiblcb = -4.953656210e-8
+ drout = 7.244550742e-01 ldrout = -3.306839609e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.121294320e-08 lalpha0 = -2.438969205e-15 walpha0 = -2.646977960e-29
+ alpha1 = 1.004650258e+00 lalpha1 = -3.109685737e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.270979414e-01 lkt1 = 7.121790080e-8
+ kt2 = 1.029101439e-03 lkt2 = -3.765776583e-8
+ at = 1.369598812e+05 lat = -5.179760850e-2
+ ute = 2.085940234e-01 lute = -1.268934703e-6
+ ua1 = 6.000602418e-09 lua1 = -4.805582324e-15 wua1 = 3.308722450e-30
+ ub1 = -4.725912025e-18 lub1 = 4.000885084e-24
+ uc1 = -7.900628978e-11 luc1 = 9.809991654e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.59 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.977095171e-01 lvth0 = -3.057139584e-9
+ k1 = 3.932297063e-01 lk1 = 8.696573668e-8
+ k2 = 5.920903785e-03 lk2 = -2.176040699e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.054929839e-01 ldsub = 5.509492874e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.573674280e-01 lvoff = 6.092439875e-9
+ nfactor = 6.240200030e-01 lnfactor = 1.201197864e-6
+ eta0 = -4.954530748e-01 leta0 = 5.033556343e-07 weta0 = -4.163336342e-23 peta0 = 1.058181320e-28
+ etab = -1.702508963e-01 letab = 8.680215367e-8
+ u0 = 2.383561950e-02 lu0 = -1.168892645e-9
+ ua = -1.286096305e-09 lua = -1.017605720e-16
+ ub = 1.987544147e-18 lub = -1.056020158e-25
+ uc = 6.258845349e-11 luc = 7.637040637e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.060478235e+04 lvsat = 6.003585447e-2
+ a0 = -5.279722970e-01 la0 = 1.035859858e-6
+ ags = 3.227856408e-01 lags = 3.945384409e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.161186290e-02 lketa = -4.252605433e-08 wketa = -1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.806822233e-01 lpclm = -1.944471501e-7
+ pdiblc1 = 5.395309339e-01 lpdiblc1 = -2.029924265e-7
+ pdiblc2 = 1.009816291e-02 lpdiblc2 = -4.337771860e-9
+ pdiblcb = -7.427084443e-02 lpdiblcb = 2.516685754e-8
+ drout = -2.184018285e-01 ldrout = 6.223425964e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.757411360e-08 lalpha0 = 1.239108811e-15
+ alpha1 = 5.406994840e-01 lalpha1 = 1.579863734e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.422128596e-01 lkt1 = -1.458275149e-8
+ kt2 = -3.610075491e-02 lkt2 = -1.274268523e-10
+ at = 1.220672433e+05 lat = -3.674433855e-2
+ ute = -8.637901776e-01 lute = -1.849837664e-7
+ ua1 = 1.402279640e-09 lua1 = -1.576620366e-16
+ ub1 = -8.575982110e-19 lub1 = 9.084763742e-26
+ uc1 = -3.564555919e-12 luc1 = 2.184446813e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.60 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.262913778e-01 lvth0 = -1.765635388e-8
+ k1 = 2.050795932e-01 lk1 = 1.830701804e-7
+ k2 = 7.863177628e-02 lk2 = -5.890010271e-08 pk2 = 1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.618143394e-01 ldsub = 7.740536886e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446112e-03 lcdscd = -1.783892580e-09 wcdscd = 6.938893904e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.109742158e-01 lvoff = -1.760456345e-8
+ nfactor = 4.519022990e+00 lnfactor = -7.883151319e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.525776721e-02 letab = -2.327665451e-08 wetab = -1.344410694e-23 petab = -1.951563910e-30
+ u0 = 2.458504396e-02 lu0 = -1.551688163e-9
+ ua = -1.881576616e-09 lua = 2.024024342e-16
+ ub = 2.589559975e-18 lub = -4.131032724e-25
+ uc = 6.187197712e-11 luc = 8.003006735e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.078372716e+04 lvsat = 2.929729196e-2
+ a0 = 1.5
+ ags = 9.337213088e-01 lags = 8.248105476e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.208158801e-02 lketa = -2.744240334e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.727091359e-01 lpclm = -1.392960087e-7
+ pdiblc1 = -8.200367215e-02 lpdiblc1 = 1.144787488e-7
+ pdiblc2 = -5.487871871e-03 lpdiblc2 = 3.623356504e-9
+ pdiblcb = 5.667376270e-02 lpdiblcb = -4.171781455e-08 ppdiblcb = 6.938893904e-30
+ drout = 1.518101815e+00 ldrout = -2.646391535e-7
+ pscbe1 = 8.089503007e+08 lpscbe1 = -4.571688292e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.876240960e-08 lalpha0 = -4.475716150e-15
+ alpha1 = 0.85
+ beta0 = 1.338015376e+01 lbeta0 = 2.450987415e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.018500067e-01 lkt1 = 1.587906831e-8
+ kt2 = -4.414385625e-02 lkt2 = 3.980876710e-9
+ at = 7.246399777e+04 lat = -1.140769520e-02 wat = -5.820766091e-17
+ ute = -1.128830784e+00 lute = -4.960473507e-8
+ ua1 = 2.259287292e-09 lua1 = -5.954095471e-16
+ ub1 = -2.127094562e-18 lub1 = 7.392886007e-25 wub1 = 7.703719778e-40
+ uc1 = -7.344148208e-11 luc1 = 5.753662374e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.61 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.364038796e-01 lvth0 = -2.029355277e-08 wvth0 = -4.358799651e-08 pvth0 = 1.136713926e-14
+ k1 = 0.90707349
+ k2 = -8.578994760e-02 lk2 = -1.602121903e-08 wk2 = -5.033029595e-08 pk2 = 1.312543656e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586434640e-01 ldsub = -3.511233284e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930381000e-02 lvoff = -2.064804189e-8
+ nfactor = -9.804248055e+00 lnfactor = 2.946993431e-06 wnfactor = 1.238450548e-05 pnfactor = -3.229705646e-12
+ eta0 = 6.941433251e-04 leta0 = -8.671466817e-16
+ etab = -0.043998
+ u0 = -4.408554454e-02 lu0 = 1.635663993e-08 wu0 = 3.886073989e-08 pu0 = -1.013433691e-14
+ ua = -7.946750893e-10 lua = -8.104626744e-17 wua = -3.912580058e-16 pua = 1.020346103e-22
+ ub = -5.749018091e-18 lub = 1.761481147e-24 wub = 5.122208891e-24 pub = -1.335800368e-30
+ uc = 3.967248006e-10 luc = -7.932192169e-17 wuc = -3.141523801e-16 puc = 8.192654260e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.010435078e+04 lvsat = 4.251376381e-02 wvsat = 8.676671606e-02 pvsat = -2.262754482e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.744150730e-01 lketa = 1.541941749e-07 wketa = 4.200474090e-07 pketa = -1.095424836e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.991951134e-01 lpclm = -4.188878082e-08 wpclm = 1.214906352e-07 ppclm = -3.168305679e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.983346087e-08 lalpha0 = 2.645242653e-14 walpha0 = 9.047174962e-14 palpha0 = -2.359376570e-20
+ alpha1 = 0.85
+ beta0 = 1.775146819e+01 lbeta0 = -8.948788635e-07 wbeta0 = -2.477202668e-06 pbeta0 = 6.460197750e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.824689802e-01 lkt1 = 6.298196792e-08 wkt1 = 2.154089277e-07 pkt1 = -5.617563261e-14
+ kt2 = -0.028878939
+ at = 1.830122700e+05 lat = -4.023713693e-02 wat = -2.154089277e-01 pat = 5.617563261e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.62 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.759269925e-01 lvth0 = -8.755409384e-09 wvth0 = -3.687103082e-08 pvth0 = 1.008563624e-14
+ k1 = 0.90707349
+ k2 = -2.991464838e-01 lk2 = 2.468422109e-08 wk2 = 1.675052933e-07 pk2 = -2.843454417e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = 3.312030375e+01 lnfactor = -5.242410110e-06 wnfactor = -3.619665670e-05 pnfactor = 6.038899963e-12
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 7.925577053e-02 lu0 = -7.175156208e-09 wu0 = -5.758045052e-08 pu0 = 8.265292041e-15
+ ua = -1.940683164e-09 lua = 1.375960290e-16 wua = 9.743342244e-16 pua = -1.585012689e-22
+ ub = 3.831602461e-18 lub = -6.636712562e-26 wub = -2.280067920e-24 pub = 7.645041575e-32
+ uc = -5.553195725e-10 luc = 1.023148161e-16 wuc = 7.330222203e-16 puc = -1.178597107e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.614499104e+05 lvsat = 2.841298718e-04 wvsat = -3.011946282e-02 pvsat = -3.272982915e-10
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 8.508406928e-01 lketa = -1.368032716e-07 wketa = -9.801106209e-07 pketa = 1.575880663e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.796361268e-01 wpclm = -4.457530670e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.132579954e-07 lalpha0 = -2.946532004e-14 walpha0 = -2.111007491e-13 palpha0 = 3.394204505e-20
+ alpha1 = 0.85
+ beta0 = 8.832221556e+00 lbeta0 = 8.067885250e-07 wbeta0 = 5.780139559e-06 pbeta0 = -9.293655192e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.153678204e-01 lkt1 = -7.015552391e-08 wkt1 = -5.026208312e-07 pkt1 = 8.081439297e-14
+ kt2 = -0.028878939
+ at = -3.956080734e+05 lat = 7.015552391e-02 wat = 5.026208312e-01 pat = -8.081439297e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.63 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.167023583e-01 lvth0 = 6.446859454e-06 wvth0 = 4.718153834e-08 pvth0 = -4.718662734e-12
+ k1 = 6.997665621e-01 lk1 = -1.317730536e-05 wk1 = -9.643851283e-08 pk1 = 9.644891469e-12
+ k2 = -7.901980754e-02 lk2 = 4.708863997e-06 wk2 = 3.446196536e-08 pk2 = -3.446568243e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.039000940e-01 lvoff = -4.378218192e-07 wvoff = -3.204212391e-09 pvoff = 3.204557998e-13
+ nfactor = 4.940526918e+00 lnfactor = -1.018436755e-04 wnfactor = -7.453460580e-07 pnfactor = 7.454264510e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.405554935e-02 lu0 = 7.949608000e-07 wu0 = 5.817944959e-09 pu0 = -5.818572482e-13
+ ua = -1.591070566e-09 lua = 5.419837178e-14 wua = 3.966524436e-16 pua = -3.966952265e-20
+ ub = 1.361072919e-18 lub = -1.127350777e-23 wub = -8.250551188e-26 pub = 8.251441093e-30
+ uc = 8.024276129e-11 luc = -3.170918107e-15 wuc = -2.320646127e-17 puc = 2.320896432e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.353357948e+00 la0 = 9.243049175e-07 wa0 = 6.764553844e-09 pa0 = -6.765283469e-13
+ ags = 3.396356791e-01 lags = 5.244886534e-07 wags = 3.838486271e-09 pags = -3.838900291e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.424943097e-08 lb0 = 1.994758229e-12 wb0 = 1.459869918e-14 pb0 = -1.460027380e-18
+ b1 = 2.963064236e-08 lb1 = -1.725750355e-12 wb1 = -1.262995682e-14 pb1 = 1.263131909e-18
+ keta = -8.748251028e-03 lketa = 4.202104218e-07 wketa = 3.075322840e-09 pketa = -3.075654544e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.606981592e-02 lpclm = 9.295484095e-06 wpclm = 6.802928501e-08 ppclm = -6.803662265e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.093461422e-03 lpdiblc2 = 3.054118263e-07 wpdiblc2 = 2.235165804e-09 ppdiblc2 = -2.235406889e-13
+ pdiblcb = 3.033677576e+00 lpdiblcb = -3.059007485e-04 wpdiblcb = -2.238743995e-06 ppdiblcb = 2.238985466e-10
+ drout = 0.56
+ pscbe1 = -5.231123437e+08 lpscbe1 = 7.481930351e+04 wpscbe1 = 5.475673639e+02 ppscbe1 = -5.476264245e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.778741884e-01 lkt1 = -8.506729023e-07 wkt1 = -6.225675686e-09 pkt1 = 6.226347188e-13
+ kt2 = -4.190194228e-02 lkt2 = 1.238534702e-06 wkt2 = 9.064254145e-09 pkt2 = -9.065231815e-13
+ at = 2.238038370e+05 lat = -4.880910095e+00 wat = -3.572109000e-02 pat = 3.572494288e-6
+ ute = -8.751456826e-01 lute = -2.402802313e-05 wute = -1.758498231e-07 pute = 1.758687902e-11
+ ua1 = 7.966636434e-10 lua1 = 3.243713395e-14 wua1 = 2.373921581e-16 pua1 = -2.374177633e-20
+ ub1 = -4.993223950e-20 lub1 = -5.195937978e-23 wub1 = -3.802663121e-25 pub1 = 3.803073276e-29
+ uc1 = 1.150093803e-10 luc1 = -8.119977561e-15 wuc1 = -5.942630444e-17 puc1 = 5.943271416e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.64 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 8.800473258e-01 lvth0 = -2.825037535e-06 wvth0 = -3.145435889e-07 pvth0 = 2.519741379e-12
+ k1 = -2.473051351e-01 lk1 = 5.774343698e-06 wk1 = 6.429234189e-07 pk1 = -5.150321923e-12
+ k2 = 2.594129521e-01 lk2 = -2.063441530e-06 wk2 = -2.297464358e-07 pk2 = 1.840449531e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.353669715e-01 lvoff = 1.918551322e-07 wvoff = 2.136141594e-08 pvoff = -1.711217318e-13
+ nfactor = -2.379123037e+00 lnfactor = 4.462827335e-05 wnfactor = 4.968973720e-06 pnfactor = -3.980538511e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.119051385e-02 lu0 = -3.483547477e-07 wu0 = -3.878629973e-08 pu0 = 3.107087468e-13
+ ua = 2.304243578e-09 lua = -2.374992594e-14 wua = -2.644349624e-15 pua = 2.118331895e-20
+ ub = 5.508298653e-19 lub = 4.940092589e-24 wub = 5.500367459e-25 pub = -4.406226663e-30
+ uc = -1.476556376e-10 luc = 1.389507982e-15 wuc = 1.547097418e-16 puc = -1.239346634e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.419789058e+00 la0 = -4.050338160e-07 wa0 = -4.509702563e-08 pa0 = 3.612626215e-13
+ ags = 3.773314254e-01 lags = -2.298328578e-07 wags = -2.558990848e-08 pags = 2.049952806e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.091166829e-07 lb0 = -8.741103958e-13 wb0 = -9.732466122e-14 pb0 = 7.796470336e-19
+ b1 = -9.440149266e-08 lb1 = 7.562301558e-13 wb1 = 8.419971215e-14 pb1 = -6.745058753e-19
+ keta = 2.145287025e-02 lketa = -1.841377530e-07 wketa = -2.050215227e-08 pketa = 1.642383543e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.920098602e-01 lpclm = -4.073315334e-06 wpclm = -4.535285667e-07 ppclm = 3.633120293e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.985692136e-02 lpdiblc2 = -1.338325861e-07 wpdiblc2 = -1.490110536e-08 ppdiblc2 = 1.193695662e-13
+ pdiblcb = -1.895184474e+01 lpdiblcb = 1.340468336e-04 wpdiblcb = 1.492495997e-05 ppdiblcb = -1.195606604e-10
+ drout = 0.56
+ pscbe1 = 4.854257521e+09 lpscbe1 = -3.278609410e+04 wpscbe1 = -3.650449093e+03 ppscbe1 = 2.924296649e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.390132610e-01 lkt1 = 3.727679960e-07 wkt1 = 4.150450457e-08 pkt1 = -3.324837042e-13
+ kt2 = 4.711331008e-02 lkt2 = -5.427304638e-07 wkt2 = -6.042836096e-08 pkt2 = 4.840786680e-13
+ at = -1.269941207e+05 lat = 2.138832764e+00 wat = 2.381406000e-01 pat = -1.907693385e-6
+ ute = -2.602073914e+00 lute = 1.052916815e-05 wute = 1.172332154e-06 pute = -9.391302005e-12
+ ua1 = 3.127966642e-09 lua1 = -1.421407145e-14 wua1 = -1.582614388e-15 pua1 = 1.267798518e-20
+ ub1 = -3.784326840e-18 lub1 = 2.276879141e-23 wub1 = 2.535108747e-24 pub1 = -2.030821366e-29
+ uc1 = -4.685849676e-10 luc1 = 3.558204046e-15 wuc1 = 3.961753629e-16 puc1 = -3.173676051e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.65 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.170743503e-01 lvth0 = 8.266129549e-8
+ k1 = 4.567336080e-01 lk1 = 1.344399904e-7
+ k2 = 1.114140034e-02 lk2 = -7.459125980e-08 wk2 = -1.734723476e-24 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.168391204e-01 lvoff = 4.343248247e-8
+ nfactor = 3.469646930e+00 lnfactor = -2.224971222e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.811640691e-02 lu0 = -3.297294898e-9
+ ua = -6.221534367e-10 lua = -3.071857119e-16
+ ub = 1.157713655e-18 lub = 7.847642182e-26
+ uc = 2.622213792e-11 luc = -3.389667350e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.501305188e+00 la0 = -1.058042092e-6
+ ags = 3.581621046e-01 lags = -7.627153156e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.285724033e-02 lketa = 9.071320047e-08 wketa = -1.734723476e-24 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.673104246e-01 lpclm = 3.611594172e-06 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.955579854e-03 lpdiblc2 = 1.560443807e-9
+ pdiblcb = -4.418017311e+00 lpdiblcb = 1.761945233e-5
+ drout = 0.56
+ pscbe1 = 7.778430133e+08 lpscbe1 = -1.308098334e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912466833e-01 lkt1 = -9.879836114e-9
+ kt2 = -2.057476356e-02 lkt2 = -4.957910604e-10
+ at = 140000.0
+ ute = -1.490445232e+00 lute = 1.624148668e-6
+ ua1 = 1.251425227e-09 lua1 = 8.185002439e-16
+ ub1 = -9.358332547e-19 lub1 = -4.988112379e-26
+ uc1 = -3.054834705e-11 luc1 = 4.918641870e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.66 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.106045433e-01 lvth0 = 1.086103068e-7
+ k1 = 4.408190516e-01 lk1 = 1.982698706e-7
+ k2 = 1.863132370e-02 lk2 = -1.046317395e-07 wk2 = 6.938893904e-24 pk2 = -1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -8.606520361e-02 lvoff = -7.999511228e-8
+ nfactor = 3.549780143e+00 lnfactor = -2.546368387e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.933554941e-02 lu0 = -8.187014548e-9
+ ua = -2.414911465e-10 lua = -1.833940696e-15
+ ub = 6.589395849e-19 lub = 2.078952480e-24
+ uc = -3.494870781e-12 luc = 1.157988951e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.515523305e+00 la0 = -1.115067914e-6
+ ags = 1.366518094e-01 lags = 8.121588595e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.846356849e-02 lketa = -7.501572108e-08 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.091009455e-01 lpclm = 9.649571892e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.381838483e-03 lpdiblc2 = 7.872383663e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.901616173e+08 lpscbe1 = 2.208614822e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957509478e-01 lkt1 = 8.185804823e-9
+ kt2 = -2.371415082e-02 lkt2 = 1.209561941e-8
+ at = 1.689553184e+05 lat = -1.161335857e-1
+ ute = -1.752105721e+00 lute = 2.673612892e-6
+ ua1 = -7.113229936e-10 lua1 = 8.690663327e-15
+ ub1 = 8.493023065e-19 lub1 = -7.209677841e-24
+ uc1 = -6.285819551e-12 luc1 = -4.812538692e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.67 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.342275017e-01 lvth0 = 6.110959292e-8
+ k1 = 6.002258295e-01 lk1 = -1.222630466e-7
+ k2 = -5.139249434e-02 lk2 = 3.617117345e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.000814656e-01 lvoff = -5.181140900e-8
+ nfactor = 2.759531280e+00 lnfactor = -9.573470380e-7
+ eta0 = 1.583042774e-01 leta0 = -1.574531447e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 2.787667965e-02 lu0 = -5.253539668e-9
+ ua = -9.177990006e-10 lua = -4.740303314e-16
+ ub = 1.500559190e-18 lub = 3.866355608e-25
+ uc = 3.787088470e-11 luc = 3.262121312e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.989214000e+04 lvsat = 2.032474338e-2
+ a0 = 1.430132279e+00 la0 = -9.433648340e-7
+ ags = 3.661307571e-01 lags = 3.507258042e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.742407017e-02 lketa = 3.736236032e-08 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.244546611e-01 lpclm = 2.667012826e-7
+ pdiblc1 = 4.418486520e-01 lpdiblc1 = -1.042565435e-7
+ pdiblc2 = 4.781655300e-03 lpdiblc2 = 1.036079606e-9
+ pdiblcb = -3.645777836e-04 lpdiblcb = -4.953656210e-8
+ drout = 7.244550742e-01 ldrout = -3.306839609e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.121294320e-08 lalpha0 = -2.438969205e-15
+ alpha1 = 1.004650258e+00 lalpha1 = -3.109685737e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.270979414e-01 lkt1 = 7.121790080e-8
+ kt2 = 1.029101439e-03 lkt2 = -3.765776583e-8
+ at = 1.369598812e+05 lat = -5.179760850e-02 wat = -1.164153218e-16
+ ute = 2.085940234e-01 lute = -1.268934703e-6
+ ua1 = 6.000602418e-09 lua1 = -4.805582324e-15
+ ub1 = -4.725912025e-18 lub1 = 4.000885084e-24 pub1 = 3.081487911e-45
+ uc1 = -7.900628978e-11 luc1 = 9.809991654e-17 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.68 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.977095171e-01 lvth0 = -3.057139584e-9
+ k1 = 3.932297063e-01 lk1 = 8.696573668e-8
+ k2 = 5.920903785e-03 lk2 = -2.176040699e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.054929839e-01 ldsub = 5.509492874e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.573674280e-01 lvoff = 6.092439875e-9
+ nfactor = 6.240200030e-01 lnfactor = 1.201197864e-6
+ eta0 = -4.954530748e-01 leta0 = 5.033556343e-07 weta0 = -1.040834086e-22 peta0 = 1.127570259e-28
+ etab = -1.702508962e-01 letab = 8.680215367e-8
+ u0 = 2.383561950e-02 lu0 = -1.168892645e-9
+ ua = -1.286096305e-09 lua = -1.017605720e-16
+ ub = 1.987544147e-18 lub = -1.056020158e-25
+ uc = 6.258845349e-11 luc = 7.637040637e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.060478235e+04 lvsat = 6.003585447e-2
+ a0 = -5.279722970e-01 la0 = 1.035859858e-6
+ ags = 3.227856408e-01 lags = 3.945384409e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.161186290e-02 lketa = -4.252605433e-08 wketa = -1.387778781e-23 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.806822233e-01 lpclm = -1.944471501e-7
+ pdiblc1 = 5.395309339e-01 lpdiblc1 = -2.029924265e-7
+ pdiblc2 = 1.009816291e-02 lpdiblc2 = -4.337771860e-9
+ pdiblcb = -7.427084443e-02 lpdiblcb = 2.516685754e-8
+ drout = -2.184018285e-01 ldrout = 6.223425964e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.757411360e-08 lalpha0 = 1.239108811e-15
+ alpha1 = 5.406994840e-01 lalpha1 = 1.579863734e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.422128596e-01 lkt1 = -1.458275149e-8
+ kt2 = -3.610075491e-02 lkt2 = -1.274268523e-10
+ at = 1.220672433e+05 lat = -3.674433855e-2
+ ute = -8.637901776e-01 lute = -1.849837664e-7
+ ua1 = 1.402279640e-09 lua1 = -1.576620366e-16
+ ub1 = -8.575982110e-19 lub1 = 9.084763742e-26
+ uc1 = -3.564555919e-12 luc1 = 2.184446813e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.69 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.262913778e-01 lvth0 = -1.765635388e-8
+ k1 = 2.050795932e-01 lk1 = 1.830701804e-7
+ k2 = 7.863177628e-02 lk2 = -5.890010271e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.618143394e-01 ldsub = 7.740536886e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446112e-03 lcdscd = -1.783892580e-09 wcdscd = 6.938893904e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.109742158e-01 lvoff = -1.760456345e-8
+ nfactor = 4.519022990e+00 lnfactor = -7.883151319e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.525776721e-02 letab = -2.327665451e-08 wetab = 4.336808690e-25 petab = -4.770489559e-30
+ u0 = 2.458504396e-02 lu0 = -1.551688163e-9
+ ua = -1.881576616e-09 lua = 2.024024342e-16
+ ub = 2.589559975e-18 lub = -4.131032724e-25
+ uc = 6.187197712e-11 luc = 8.003006735e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.078372716e+04 lvsat = 2.929729196e-2
+ a0 = 1.5
+ ags = 9.337213088e-01 lags = 8.248105476e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.208158801e-02 lketa = -2.744240334e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.727091359e-01 lpclm = -1.392960087e-7
+ pdiblc1 = -8.200367215e-02 lpdiblc1 = 1.144787488e-7
+ pdiblc2 = -5.487871871e-03 lpdiblc2 = 3.623356504e-09 wpdiblc2 = 1.734723476e-24 ppdiblc2 = 8.673617380e-31
+ pdiblcb = 5.667376270e-02 lpdiblcb = -4.171781455e-08 ppdiblcb = 6.938893904e-30
+ drout = 1.518101815e+00 ldrout = -2.646391535e-7
+ pscbe1 = 8.089503007e+08 lpscbe1 = -4.571688292e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.876240960e-08 lalpha0 = -4.475716150e-15
+ alpha1 = 0.85
+ beta0 = 1.338015376e+01 lbeta0 = 2.450987415e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.018500067e-01 lkt1 = 1.587906831e-8
+ kt2 = -4.414385625e-02 lkt2 = 3.980876710e-9
+ at = 7.246399777e+04 lat = -1.140769520e-2
+ ute = -1.128830784e+00 lute = -4.960473507e-8
+ ua1 = 2.259287292e-09 lua1 = -5.954095471e-16
+ ub1 = -2.127094562e-18 lub1 = 7.392886007e-25 pub1 = 1.925929944e-46
+ uc1 = -7.344148208e-11 luc1 = 5.753662374e-17 puc1 = 1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.70 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.875346872e-01 lvth0 = -7.549151562e-9
+ k1 = 0.90707349
+ k2 = -1.422183479e-01 lk2 = -1.305482221e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586434640e-01 ldsub = -3.511233285e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930381000e-02 lvoff = -2.064804189e-8
+ nfactor = 4.080785197e+00 lnfactor = -6.740288509e-7
+ eta0 = 6.941433251e-04 leta0 = -8.671466817e-16
+ etab = -0.043998
+ u0 = -5.163712314e-04 lu0 = 4.994409498e-9
+ ua = -1.233338581e-09 lua = 3.335102999e-17
+ ub = -6.193647714e-21 lub = 2.638329318e-25
+ uc = 4.450918314e-11 luc = 1.253098032e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.373838699e+05 lvsat = 1.714462714e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.034740047e-01 lketa = 3.137933746e-08 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.354057609e-01 lpclm = -7.741061073e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.16e-8
+ alpha1 = 0.85
+ beta0 = 1.497412343e+01 lbeta0 = -1.705862324e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.24096074
+ kt2 = -0.028878939
+ at = -5.849597014e+04 lat = 2.274483099e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.71 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 7.299937748e-01 lvth0 = -3.472835104e-08 wvth0 = -1.742881241e-07 pvth0 = 3.325173404e-14
+ k1 = 0.90707349
+ k2 = 1.769009749e-02 lk2 = -3.181377489e-08 wk2 = -1.150913923e-07 pk2 = 2.195782638e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587461769e-01 ldsub = -2.310740521e-11 wdsub = -1.080280217e-10 pdsub = 2.061023415e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = -6.481886456e+00 lnfactor = 1.341181023e-06 wnfactor = -8.741959909e-07 pnfactor = 1.667843563e-13
+ eta0 = -1.632446765e-02 leta0 = 3.246912159e-09 weta0 = 1.517944113e-08 peta0 = -2.896024855e-15
+ etab = -0.043998
+ u0 = 3.603765658e-02 lu0 = -1.979587253e-09 wu0 = -1.903283172e-08 pu0 = 3.631197832e-15
+ ua = -2.620746877e-09 lua = 2.980491091e-16 wua = 1.580904812e-15 pua = -3.016145055e-22
+ ub = 1.618074477e-17 lub = -2.824408301e-24 wub = -1.329466311e-23 pub = 2.536435597e-30
+ uc = 1.680052029e-10 luc = -1.103033130e-17 wuc = 8.786570671e-17 puc = -1.676354672e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.896559766e+05 lvsat = -1.263783590e-01 wvsat = -5.904365558e-01 pvsat = 1.126470287e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.635612593e-06 lb0 = 1.075195984e-12 wb0 = 5.026583212e-12 pb0 = -9.590017046e-19
+ b1 = 3.860048929e-06 lb1 = -7.364432949e-13 wb1 = -3.442901161e-12 pb1 = 6.568573409e-19
+ keta = -9.099966544e-01 lketa = 1.661739677e-07 wketa = 5.904365558e-07 pketa = -1.126470287e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.092221223e-02 lpclm = 7.390627578e-09 wpclm = 3.455147252e-08 ppclm = -6.591937237e-15
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.342008000e-08 lalpha0 = 8.589200983e-15
+ alpha1 = 0.85
+ beta0 = 2.021621011e+01 lbeta0 = -1.170702981e-06 wbeta0 = -4.373604117e-06 pbeta0 = 8.344224351e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.385031506e-01 lkt1 = 1.140027264e-07 wkt1 = 4.373604117e-07 pkt1 = -8.344224351e-14
+ kt2 = -0.028878939
+ at = 4.866397872e+05 lat = -8.125943962e-02 wat = -2.842842676e-01 pat = 5.423745828e-8
+ ute = -9.316384008e-02 lute = -2.338806196e-07 wute = -1.093401029e-06 pute = 2.086056088e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.72 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.73 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.503030477e-01 lvth0 = 6.175519114e-7
+ k1 = 6.310871457e-01 lk1 = -1.262268888e-6
+ k2 = -5.447745820e-02 lk2 = 4.510673736e-07 wk2 = -2.775557562e-23 pk2 = 2.220446049e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.061819981e-01 lvoff = -4.193944404e-8
+ nfactor = 4.409723085e+00 lnfactor = -9.755720117e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.819884287e-02 lu0 = 7.615018832e-8
+ ua = -1.308591527e-09 lua = 5.191722935e-15
+ ub = 1.302315995e-18 lub = -1.079901978e-24
+ uc = 6.371610434e-11 luc = -3.037458086e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.358175376e+00 la0 = 8.854020668e-8
+ ags = 3.423692862e-01 lags = 5.024135747e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.385285691e-08 lb0 = 1.910801322e-13
+ b1 = 2.063612306e-08 lb1 = -1.653115657e-13
+ keta = -6.558136603e-03 lketa = 4.025242849e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.762224597e-02 lpclm = 8.904248667e-07 ppclm = 2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -5.016711857e-04 lpdiblc2 = 2.925574203e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = 1.439339104e+00 lpdiblcb = -2.930257643e-05 wpdiblcb = -2.498001805e-22 ppdiblcb = -5.329070518e-27
+ drout = 0.56
+ pscbe1 = -1.331581032e+08 lpscbe1 = 7.167025156e+03 ppscbe1 = 1.907348633e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.823078504e-01 lkt1 = -8.148691321e-8
+ kt2 = -3.544676512e-02 lkt2 = 1.186406308e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.000378464e+00 lute = -2.301671335e-6
+ ua1 = 9.657242647e-10 lua1 = 3.107189510e-15
+ ub1 = -3.207417704e-19 lub1 = -4.977247376e-24
+ uc1 = 7.268848809e-11 luc1 = -7.778217749e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.74 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.170743503e-01 lvth0 = 8.266129549e-8
+ k1 = 4.567336080e-01 lk1 = 1.344399904e-7
+ k2 = 1.114140034e-02 lk2 = -7.459125980e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.168391204e-01 lvoff = 4.343248247e-8
+ nfactor = 3.469646930e+00 lnfactor = -2.224971222e-06 wnfactor = -3.552713679e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.811640691e-02 lu0 = -3.297294898e-9
+ ua = -6.221534367e-10 lua = -3.071857119e-16
+ ub = 1.157713655e-18 lub = 7.847642182e-26
+ uc = 2.622213792e-11 luc = -3.389667350e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.501305188e+00 la0 = -1.058042092e-6
+ ags = 3.581621046e-01 lags = -7.627153156e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.285724033e-02 lketa = 9.071320047e-08 wketa = -3.469446952e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.673104246e-01 lpclm = 3.611594172e-06 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.955579854e-03 lpdiblc2 = 1.560443807e-9
+ pdiblcb = -4.418017311e+00 lpdiblcb = 1.761945233e-5
+ drout = 0.56
+ pscbe1 = 7.778430133e+08 lpscbe1 = -1.308098334e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912466833e-01 lkt1 = -9.879836114e-9
+ kt2 = -2.057476356e-02 lkt2 = -4.957910604e-10
+ at = 140000.0
+ ute = -1.490445232e+00 lute = 1.624148668e-6
+ ua1 = 1.251425227e-09 lua1 = 8.185002439e-16
+ ub1 = -9.358332547e-19 lub1 = -4.988112379e-26
+ uc1 = -3.054834705e-11 luc1 = 4.918641870e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.75 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.106045433e-01 lvth0 = 1.086103068e-7
+ k1 = 4.408190516e-01 lk1 = 1.982698706e-7
+ k2 = 1.863132370e-02 lk2 = -1.046317395e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -8.606520361e-02 lvoff = -7.999511228e-8
+ nfactor = 3.549780143e+00 lnfactor = -2.546368387e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.933554941e-02 lu0 = -8.187014548e-9
+ ua = -2.414911465e-10 lua = -1.833940696e-15
+ ub = 6.589395849e-19 lub = 2.078952480e-24
+ uc = -3.494870781e-12 luc = 1.157988951e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.515523305e+00 la0 = -1.115067914e-6
+ ags = 1.366518094e-01 lags = 8.121588595e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.846356849e-02 lketa = -7.501572108e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.091009455e-01 lpclm = 9.649571892e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.381838483e-03 lpdiblc2 = 7.872383663e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.901616173e+08 lpscbe1 = 2.208614822e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957509478e-01 lkt1 = 8.185804823e-9
+ kt2 = -2.371415082e-02 lkt2 = 1.209561941e-8
+ at = 1.689553184e+05 lat = -1.161335857e-1
+ ute = -1.752105721e+00 lute = 2.673612892e-6
+ ua1 = -7.113229936e-10 lua1 = 8.690663327e-15
+ ub1 = 8.493023065e-19 lub1 = -7.209677841e-24 pub1 = -3.081487911e-45
+ uc1 = -6.285819551e-12 luc1 = -4.812538692e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.76 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.342275017e-01 lvth0 = 6.110959292e-8
+ k1 = 6.002258295e-01 lk1 = -1.222630466e-7
+ k2 = -5.139249434e-02 lk2 = 3.617117345e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.000814656e-01 lvoff = -5.181140900e-8
+ nfactor = 2.759531280e+00 lnfactor = -9.573470380e-7
+ eta0 = 1.583042774e-01 leta0 = -1.574531447e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 2.787667965e-02 lu0 = -5.253539668e-9
+ ua = -9.177990006e-10 lua = -4.740303314e-16
+ ub = 1.500559190e-18 lub = 3.866355608e-25
+ uc = 3.787088470e-11 luc = 3.262121312e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.989214000e+04 lvsat = 2.032474338e-2
+ a0 = 1.430132279e+00 la0 = -9.433648340e-7
+ ags = 3.661307571e-01 lags = 3.507258042e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.742407017e-02 lketa = 3.736236032e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.244546611e-01 lpclm = 2.667012826e-7
+ pdiblc1 = 4.418486520e-01 lpdiblc1 = -1.042565435e-07 wpdiblc1 = 4.440892099e-22
+ pdiblc2 = 4.781655300e-03 lpdiblc2 = 1.036079606e-9
+ pdiblcb = -3.645777836e-04 lpdiblcb = -4.953656210e-8
+ drout = 7.244550742e-01 ldrout = -3.306839609e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.121294320e-08 lalpha0 = -2.438969205e-15
+ alpha1 = 1.004650258e+00 lalpha1 = -3.109685737e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.270979414e-01 lkt1 = 7.121790080e-8
+ kt2 = 1.029101439e-03 lkt2 = -3.765776583e-8
+ at = 1.369598812e+05 lat = -5.179760850e-02 wat = 1.164153218e-16
+ ute = 2.085940234e-01 lute = -1.268934703e-6
+ ua1 = 6.000602418e-09 lua1 = -4.805582324e-15
+ ub1 = -4.725912025e-18 lub1 = 4.000885084e-24 pub1 = -3.081487911e-45
+ uc1 = -7.900628978e-11 luc1 = 9.809991654e-17 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.77 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.236711974e-01 lvth0 = -2.929884253e-08 wvth0 = -1.900218456e-08 pvth0 = 1.920714212e-14
+ k1 = -1.781222905e-01 lk1 = 6.644803362e-07 wk1 = 4.181908098e-07 pk1 = -4.227014158e-13
+ k2 = 1.938136854e-01 lk2 = -2.116798002e-07 wk2 = -1.375247395e-07 pk2 = 1.390080813e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.858104465e-01 ldsub = 7.498976201e-08 wdsub = 1.440627898e-08 pdsub = -1.456166511e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.457251973e-01 lvoff = -5.675363950e-09 wvoff = -8.521321219e-09 pvoff = 8.613232189e-15
+ nfactor = -4.413252793e-01 lnfactor = 2.278033960e-06 wnfactor = 7.797603032e-07 pnfactor = -7.881707978e-13
+ eta0 = -4.954530747e-01 leta0 = 5.033556341e-07 weta0 = -9.483244051e-17 peta0 = 9.585536531e-23
+ etab = -1.722682838e-01 letab = 8.884130080e-08 wetab = 1.476590533e-09 petab = -1.492517039e-15
+ u0 = 4.889606133e-03 lu0 = 1.798147243e-08 wu0 = 1.386719346e-08 pu0 = -1.401676501e-14
+ ua = -1.982656674e-09 lua = 6.023128972e-16 wua = 5.098348240e-16 pua = -5.153339024e-22
+ ub = 1.028495504e-18 lub = 8.637909260e-25 wub = 7.019583914e-25 pub = -7.095297147e-31
+ uc = -9.882192274e-11 luc = 1.707883892e-16 wuc = 1.181414195e-16 puc = -1.194156928e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.562863936e+06 lvsat = -1.488750246e+00 wvsat = -1.121509507e+00 pvsat = 1.133606108e-6
+ a0 = -1.272953194e+00 la0 = 1.788876119e-06 wa0 = 5.452753582e-07 pa0 = -5.511566982e-13
+ ags = -5.738737879e+00 lags = 6.521441554e-06 wags = 4.436623033e-06 pags = -4.484476449e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.480044889e-17 lb0 = 1.496008653e-23 wb0 = 1.083292215e-23 pb0 = -1.094976605e-29
+ b1 = -8.560766018e-17 lb1 = 8.653102440e-23 wb1 = 6.265898593e-23 pb1 = -6.333482575e-29
+ keta = 2.099747374e-01 lketa = -2.025970308e-07 wketa = -1.159108555e-07 pketa = 1.171610700e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.695849122e-01 lpclm = 1.200056566e-07 wpclm = 2.277020771e-07 ppclm = -2.301580717e-13
+ pdiblc1 = -1.646971660e-01 lpdiblc1 = 5.088314777e-07 wpdiblc1 = 5.154470816e-07 ppdiblc1 = -5.210066939e-13
+ pdiblc2 = 3.137653477e-05 lpdiblc2 = 5.837594878e-09 wpdiblc2 = 7.368203088e-09 ppdiblc2 = -7.447676527e-15
+ pdiblcb = -5.236170481e-01 lpdiblcb = 4.793597093e-07 wpdiblcb = 3.288908655e-07 ppdiblcb = -3.324382824e-13
+ drout = -2.184024743e-01 ldrout = 6.223432491e-07 wdrout = 4.726609921e-13 pdrout = -4.777591138e-19
+ pscbe1 = -1.543739537e+09 lpscbe1 = 2.369019111e+03 wpscbe1 = 1.715457967e+03 ppscbe1 = -1.733960896e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.501090235e-05 lalpha0 = -2.525155931e-11 walpha0 = -1.828609740e-11 palpha0 = 1.848333125e-17
+ alpha1 = 5.406994840e-01 lalpha1 = 1.579863734e-7
+ beta0 = 4.070255265e+01 lbeta0 = -2.713207642e-05 wbeta0 = -1.964692325e-05 pbeta0 = 1.985883496e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.950657684e-01 lkt1 = 3.884022869e-08 wkt1 = 3.868473517e-08 pkt1 = -3.910198873e-14
+ kt2 = -3.847883851e-02 lkt2 = 2.276306765e-09 wkt2 = 1.740595491e-09 pkt2 = -1.759369554e-15
+ at = -1.327699865e+05 lat = 2.208415655e-01 wat = 1.865235232e-01 pat = -1.885353659e-7
+ ute = -1.408217571e+00 lute = 3.653158208e-07 wute = 3.984838308e-07 pute = -4.027818774e-13
+ ua1 = -2.887400415e-10 lua1 = 1.551596983e-15 wua1 = 1.237711418e-15 pua1 = -1.251061373e-21
+ ub1 = -5.486267437e-19 lub1 = -2.214563962e-25 wub1 = -2.261461040e-25 pub1 = 2.285853159e-31
+ uc1 = -2.195792942e-10 luc1 = 2.401891414e-16 wuc1 = 1.581080994e-16 puc1 = -1.598134534e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.78 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.551590434e-01 lvth0 = 5.696206559e-09 wvth0 = 5.206403179e-08 pvth0 = -1.709248626e-14
+ k1 = 1.347783586e+00 lk1 = -1.149310229e-07 wk1 = -8.363816188e-07 pk1 = 2.181166167e-13
+ k2 = -2.966823963e-01 lk2 = 3.885873141e-08 wk2 = 2.747044530e-07 pk2 = -7.155281897e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.011794144e-01 ldsub = 6.713950838e-08 wdsub = -2.881255807e-08 pdsub = 7.513911793e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446104e-03 lcdscd = -1.783892576e-09 wcdscd = 5.922227986e-18 pcdscd = -3.024993450e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.342586770e-01 lvoff = -1.153230201e-08 wvoff = 1.704264226e-08 pvoff = -4.444482458e-15
+ nfactor = 6.649713556e+00 lnfactor = -1.343969402e-06 wnfactor = -1.559520608e-06 pnfactor = 4.067011416e-13
+ eta0 = 1.000416472e+00 leta0 = -2.607135882e-07 weta0 = -7.090861232e-17 peta0 = 8.363554294e-23
+ etab = 4.929254235e-02 letab = -2.432886737e-08 wetab = -2.953181039e-09 petab = 7.701482633e-16
+ u0 = 7.336237544e-02 lu0 = -1.699345951e-08 wu0 = -3.570168978e-08 pu0 = 1.130232659e-14
+ ua = -4.884558750e-10 lua = -1.609039523e-16 wua = -1.019669650e-15 pua = 2.659155701e-22
+ ub = 4.507657262e-18 lub = -9.133161921e-25 wub = -1.403916784e-24 pub = 3.661218427e-31
+ uc = 3.846927297e-10 luc = -7.618412607e-17 wuc = -2.362828391e-16 puc = 6.161925649e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.515487836e+06 lvsat = 5.944147421e-01 wvsat = 1.907613558e+00 pvsat = -4.136275455e-7
+ a0 = 2.989961792e+00 la0 = -3.885611752e-07 wa0 = -1.090550714e-06 pa0 = 2.844003581e-13
+ ags = 1.305676835e+01 lags = -3.079039890e-06 wags = -8.873246066e-06 pags = 2.314018348e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.960089777e-17 lb0 = -7.719499726e-24 wb0 = -2.166584431e-23 pb0 = 5.650148874e-30
+ b1 = 1.712153204e-16 lb1 = -4.465055854e-23 wb1 = -1.253179719e-22 pb1 = 3.268117261e-29
+ keta = -2.946441610e-01 lketa = 5.515523782e-08 wketa = 2.318217109e-07 pketa = -6.045585669e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.394903759e+00 lpclm = -3.015556556e-07 wpclm = -4.554041545e-07 ppclm = 1.187630279e-13
+ pdiblc1 = 1.326452528e+00 lpdiblc1 = -2.528269100e-07 wpdiblc1 = -1.030894164e-06 ppdiblc1 = 2.688427654e-13
+ pdiblc2 = 1.464570088e-02 lpdiblc2 = -1.627197395e-09 wpdiblc2 = -1.473640617e-08 ppdiblc2 = 3.843048417e-15
+ pdiblcb = 9.553661700e-01 lpdiblcb = -2.760842127e-07 wpdiblcb = -6.577817310e-07 ppdiblcb = 1.715402665e-13
+ drout = 1.518103104e+00 ldrout = -2.646394890e-07 wdrout = -9.435148982e-13 pdrout = 2.456037045e-19
+ pscbe1 = 5.496429374e+09 lpscbe1 = -1.227000606e+03 wpscbe1 = -3.430915933e+03 ppscbe1 = 8.947348424e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -4.992789407e-05 lalpha0 = 1.302612876e-11 walpha0 = 3.657219481e-11 palpha0 = -9.537516395e-18
+ alpha1 = 0.85
+ beta0 = -4.030495154e+01 lbeta0 = 1.424542261e-05 wbeta0 = 3.929384649e-05 pbeta0 = -1.024728505e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.961441894e-01 lkt1 = -1.168752896e-08 wkt1 = -7.736947029e-08 pkt1 = 2.017687467e-14
+ kt2 = -3.938768905e-02 lkt2 = 2.740534894e-09 wkt2 = -3.481190971e-09 pkt2 = 9.078458658e-16
+ at = 5.821384572e+05 lat = -1.443236588e-01 wat = -3.730470465e-01 pat = 9.728544706e-8
+ ute = -3.997599746e-02 lute = -3.335628195e-07 wute = -7.969676618e-07 pute = 2.078380087e-13
+ ua1 = 5.641326653e-09 lua1 = -1.477398063e-15 wua1 = -2.475422833e-15 pua1 = 6.455556185e-22
+ ub1 = -2.745037501e-18 lub1 = 9.004394689e-25 wub1 = 4.522922110e-25 pub1 = -1.179514773e-31
+ uc1 = 3.585879945e-10 luc1 = -5.513061536e-17 wuc1 = -3.162161989e-16 puc1 = 8.246475765e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.79 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 1.197330485e+00 lvth0 = -1.617731150e-07 wvth0 = -4.463290577e-07 pvth0 = 1.128814540e-13
+ k1 = 9.070734932e-01 lk1 = -6.073390679e-16 wk1 = -2.329997528e-15 pk1 = 4.445310786e-22
+ k2 = -6.408110130e-02 lk2 = -2.180042990e-08 wk2 = -5.719115118e-08 pk2 = 1.500090805e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587285471e-01 ldsub = -2.569974795e-11 wdsub = -6.227504236e-11 pdsub = 1.624048392e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000032e-03 lcdscd = -6.426701185e-18 wcdscd = -2.371471769e-17 pcdscd = 4.703908270e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930381134e-02 lvoff = -2.064804160e-08 wvoff = 9.804734802e-16 pvoff = -2.105716712e-22
+ nfactor = 2.776520619e+01 lnfactor = -6.850594264e-06 wnfactor = -1.733538563e-05 pnfactor = 4.520825876e-12
+ eta0 = -1.126128123e-02 leta0 = 3.117806392e-09 weta0 = 8.750557806e-09 peta0 = -2.282022903e-15
+ etab = -4.399799986e-02 letab = -2.622341233e-17 wetab = -1.006036365e-16 petab = 1.919375769e-23
+ u0 = -3.519381827e-02 lu0 = 1.131647602e-08 wu0 = 2.538153316e-08 pu0 = -4.627322791e-15
+ ua = -1.822370922e-09 lua = 1.869624172e-16 wua = 4.311316193e-16 pua = -1.124330899e-22
+ ub = 8.025675296e-19 lub = 5.291933898e-26 wub = -5.919581861e-25 pub = 1.543744078e-31
+ uc = -5.270664684e-10 luc = 1.615899082e-16 wuc = 4.183545098e-16 puc = -1.091009992e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.200529879e+05 lvsat = 4.795466975e-02 wvsat = 4.080058742e-01 pvsat = -2.255085611e-8
+ a0 = 1.500000010e+00 la0 = -1.855308795e-15 wa0 = -7.117712642e-15 pa0 = 1.357959967e-21
+ ags = 1.250000002e+00 lags = -3.972386864e-16 wags = -1.523968507e-15 pags = 2.907523111e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.673484566e-07 lb0 = 6.972073460e-14 wb0 = 1.956808905e-13 pb0 = -5.103083672e-20
+ b1 = 1.831174339e-07 lb1 = -4.775446311e-14 wb1 = -1.340295096e-13 pb1 = 3.495301970e-20
+ keta = 3.206758066e-03 lketa = -2.252011195e-08 wketa = -1.512762640e-07 pketa = 3.945073181e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.389742803e+00 lpclm = -3.002097506e-07 wpclm = -6.253166196e-07 ppclm = 1.630738200e-13
+ pdiblc1 = 3.569721483e-01 lpdiblc1 = 3.176248153e-16 wpdiblc1 = 1.218537271e-15 ppdiblc1 = -2.324798132e-22
+ pdiblc2 = 8.406112145e-03 lpdiblc2 = -8.516243266e-18 wpdiblc2 = -3.267175419e-17 ppdiblc2 = 6.233315947e-24
+ pdiblcb = -1.032957699e-01 lpdiblcb = -2.521605147e-17 wpdiblcb = -9.673883916e-17 ppdiblcb = 1.845640307e-23
+ drout = 5.033266688e-01 ldrout = -1.682273876e-15 wdrout = -6.453880985e-15 pdrout = 1.231310165e-21
+ pscbe1 = 7.914198809e+08 lpscbe1 = -1.661944389e-07 wpscbe1 = -6.375885010e-07 ppscbe1 = 1.216430664e-13
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.662765292e-07 lalpha0 = -3.772961370e-14 walpha0 = -1.058933814e-13 palpha0 = 2.761551162e-20
+ alpha1 = 0.85
+ beta0 = 1.123895178e+01 lbeta0 = 8.034942409e-07 wbeta0 = 2.733891654e-06 pbeta0 = -7.129606690e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.003724933e-02 lkt1 = -4.196659342e-08 wkt1 = -1.177850524e-07 pkt1 = 3.071669265e-14
+ kt2 = -2.887893895e-02 lkt2 = -1.008054751e-17 wkt2 = -3.867306475e-17 pkt2 = 7.378278544e-24
+ at = -1.790597490e+05 lat = 5.418617662e-02 wat = 8.824448777e-02 pat = -2.301292699e-8
+ ute = -1.262490799e+00 lute = -1.474807435e-08 wute = -4.139251161e-08 pute = 1.079458756e-14
+ ua1 = -2.384732603e-11 lua1 = -1.902030267e-24 wua1 = -7.296954800e-24 pua1 = 1.392156823e-30
+ ub1 = 7.077531842e-19 lub1 = -2.701925638e-33 wub1 = -1.036567544e-32 pub1 = 1.977626141e-39
+ uc1 = 1.471862498e-10 luc1 = 3.912212746e-26 wuc1 = 1.500877862e-25 puc1 = -2.863471806e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.80 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = -7.924619035e-01 lvth0 = 2.178514156e-07 wvth0 = 9.400459055e-07 pvth0 = -1.516194797e-13
+ k1 = 0.90707349
+ k2 = -4.083638064e-01 lk2 = 4.388389027e-08 wk2 = 1.967510936e-07 pk2 = -3.344771707e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584000555e-01 ldsub = 3.697184834e-11 wdsub = 1.453092562e-10 pdsub = -2.336369407e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999992e-03 lcdscd = 1.230168745e-18 wcdscd = 5.660125146e-18 pcdscd = -9.003995466e-25
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075299989e-01 lvoff = -1.721580656e-16 wvoff = -7.836993277e-16 pvoff = 1.260079818e-22
+ nfactor = -6.537596072e+01 lnfactor = 1.091943640e-05 wnfactor = 4.223226157e-05 pnfactor = -6.843847262e-12
+ eta0 = 3.231038961e-02 leta0 = -5.195057784e-09 weta0 = -2.041796604e-08 peta0 = 3.282923088e-15
+ etab = -0.043998
+ u0 = -2.740290011e-02 lu0 = 9.830077904e-09 wu0 = 2.740134182e-08 pu0 = -5.012674006e-15
+ ua = 2.095541840e-09 lua = -5.605204870e-16 wua = -1.871097821e-15 pua = 3.268000561e-22
+ ub = -1.273520232e-17 lub = 2.635736298e-24 wub = 7.869843871e-24 pub = -1.460018959e-30
+ uc = 1.621727993e-09 luc = -2.483699919e-16 wuc = -9.761605222e-16 puc = 1.569529457e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.655766123e+06 lvsat = 4.744974360e-01 wvsat = 2.004571333e+00 pvsat = -3.271531937e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.132305965e-06 lb0 = -9.604577340e-13 wb0 = -2.854800955e-12 pb0 = 5.309583927e-19
+ b1 = -3.515314392e-06 lb1 = 6.578545512e-13 wb1 = 1.955363265e-12 pb1 = -3.636738702e-19
+ keta = -5.855695136e-01 lketa = 8.981015782e-08 wketa = 3.529779498e-07 pketa = -5.675391264e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.072893516e+00 lpclm = 1.696267822e-07 wpclm = 8.863854464e-07 ppclm = -1.253377703e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.609986601e-07 lalpha0 = 6.286711056e-14 walpha0 = 2.470845653e-13 palpha0 = -3.972773891e-20
+ alpha1 = 0.85
+ beta0 = 2.005574672e+01 lbeta0 = -8.786267981e-07 wbeta0 = -4.256155829e-06 pbeta0 = 6.206425301e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.739035193e-01 lkt1 = 3.317757676e-08 wkt1 = 1.704982743e-07 pkt1 = -2.428373011e-14
+ kt2 = -0.028878939
+ at = 3.795527042e+05 lat = -5.238925888e-02 wat = -2.059038048e-01 pat = 3.310644915e-8
+ ute = -2.444085418e+00 lute = 2.106836366e-07 wute = 6.273137034e-07 pute = -1.167851964e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.81 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.82 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.225219353e-01 lvth0 = 1.173473807e-06 wvth0 = 1.755577392e-08 pvth0 = -3.513048351e-13
+ k1 = 7.428610218e-01 lk1 = -3.498952003e-06 wk1 = -7.063348909e-08 pk1 = 1.413431635e-12
+ k2 = -1.089747373e-01 lk2 = 1.541600763e-06 wk2 = 3.443857457e-08 pk2 = -6.891429458e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.334255931e-01 lvoff = 5.032263052e-07 wvoff = 1.721609947e-08 pvoff = -3.445076822e-13
+ nfactor = 4.723261510e+00 lnfactor = -1.602987046e-05 wnfactor = -1.981349644e-07 pnfactor = 3.964836372e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.021888796e-02 lu0 = 2.358353582e-07 wu0 = 5.042788863e-09 pu0 = -1.009101688e-13
+ ua = -1.738043863e-09 lua = 1.378540172e-14 wua = 2.713846733e-16 pua = -5.430620621e-21
+ ub = 1.361365732e-18 lub = -2.261533625e-24 wub = -3.731541830e-26 pub = 7.467108501e-31
+ uc = 6.580234079e-11 luc = -3.454930397e-16 wuc = -1.318359571e-18 puc = 2.638141124e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.160292432e+00 la0 = 4.048333449e-06 wa0 = 1.250485645e-07 pa0 = -2.502320063e-12
+ ags = 4.724837131e-01 lags = -2.553450595e-06 wags = -8.222347004e-08 pags = 1.645356263e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.630435158e-08 lb0 = 1.640891487e-12 wb0 = 4.578441793e-14 pb0 = -9.161821893e-19
+ b1 = 4.155395972e-08 lb1 = -5.838939187e-13 wb1 = -1.321865036e-14 pb1 = 2.645155835e-19
+ keta = -3.007770829e-02 lketa = 5.108975443e-07 wketa = 1.486276997e-08 pketa = -2.974157093e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.347719931e-01 lpclm = 3.034575526e-06 wpclm = 6.771135399e-08 ppclm = -1.354957415e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -6.833560397e-03 lpdiblc2 = 1.559618220e-07 wpdiblc2 = 4.001323413e-09 ppdiblc2 = -8.006962654e-14
+ pdiblcb = 1.025680820e+01 lpdiblcb = -2.057470637e-04 wpdiblcb = -5.572040884e-06 ppdiblcb = 1.115009177e-10
+ drout = 0.56
+ pscbe1 = -4.809228255e+08 lpscbe1 = 1.412607059e+04 wpscbe1 = 2.197636565e+02 ppscbe1 = -4.397643502e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.769214211e-01 lkt1 = -1.892735985e-07 wkt1 = -3.403857081e-09 pkt1 = 6.811385562e-14
+ kt2 = -3.518413649e-02 lkt2 = 1.133852255e-07 wkt2 = -1.659634346e-10 pkt2 = 3.321058774e-15
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -9.095327154e-01 lute = -4.119566177e-06 wute = -5.740833584e-08 pute = 1.148785923e-12
+ ua1 = 5.818406794e-10 lua1 = 1.078900178e-14 wua1 = 2.425883218e-16 pua1 = -4.854382994e-21
+ ub1 = 4.726390747e-20 lub1 = -1.234133024e-23 wub1 = -2.325545640e-25 pub1 = 4.653599614e-30
+ uc1 = 9.210253818e-11 luc1 = -1.166312177e-15 wuc1 = -1.226835950e-17 puc1 = 2.454995166e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.83 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.011796457e-01 lvth0 = -2.577148786e-07 wvth0 = -5.314882753e-08 pvth0 = 2.150945964e-13
+ k1 = 5.792489871e-01 lk1 = -2.188291007e-06 wk1 = -7.742138855e-08 pk1 = 1.467808045e-12
+ k2 = -4.773521515e-02 lk2 = 1.051024056e-06 wk2 = 3.720601738e-08 pk2 = -7.113123380e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.098697167e-01 lvoff = 3.145252203e-07 wvoff = -4.404189257e-09 pvoff = -1.713121760e-13
+ nfactor = 3.087241344e-01 lnfactor = 1.933404375e-05 wnfactor = 1.997488264e-06 pnfactor = -1.362383145e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.463195597e-02 lu0 = -1.199482252e-07 wu0 = -1.675602394e-08 pu0 = 7.371545566e-14
+ ua = 1.499634463e-09 lua = -1.215094648e-14 wua = -1.340825671e-15 pua = 7.484451432e-21
+ ub = -1.239628140e-20 lub = 8.743379878e-24 wub = 7.394299124e-25 pub = -5.475629771e-30
+ uc = 1.271930437e-10 luc = -8.372808228e-16 wuc = -6.380674640e-17 puc = 5.269625056e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.049635017e+00 la0 = -3.075999680e-06 wa0 = -3.465071653e-07 pa0 = 1.275211975e-12
+ ags = 3.423043678e-01 lags = -1.510611718e-06 wags = 1.002101137e-08 pags = 9.064054629e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.785793739e-09 lb0 = 8.070476086e-13 wb0 = -4.920092209e-15 pb0 = -5.099992094e-19
+ b1 = -3.667485703e-08 lb1 = 4.278039133e-14 wb1 = 2.317601575e-14 pb1 = -2.703429826e-20
+ keta = 1.541054804e-02 lketa = 1.465008573e-07 wketa = -1.786332004e-08 pketa = -3.525400558e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.642642992e+00 lpclm = -1.120391555e-05 wpclm = -1.270153882e-06 ppclm = 9.362394691e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.081681516e-02 lpdiblc2 = -1.456472794e-07 wpdiblc2 = -1.760640615e-08 ppdiblc2 = 9.302527093e-14
+ pdiblcb = -3.087042461e+01 lpdiblcb = 1.237143972e-04 wpdiblcb = 1.671612265e-05 ppdiblcb = -6.704479071e-11
+ drout = 0.56
+ pscbe1 = 1.615700996e+09 lpscbe1 = -2.669534166e+03 wpscbe1 = -5.294692710e+02 ppscbe1 = 1.604301145e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.214738207e-01 lkt1 = 1.676261404e-07 wkt1 = 1.910149537e-08 pkt1 = -1.121717067e-13
+ kt2 = -8.604929512e-02 lkt2 = 5.208551261e-07 wkt2 = 4.137545168e-08 pkt2 = -3.294583278e-13
+ at = 140000.0
+ ute = -3.054447269e+00 lute = 1.306288530e-05 wute = 9.883429350e-07 pute = -7.228503717e-12
+ ua1 = -3.546451147e-10 lua1 = 1.829098907e-14 wua1 = 1.014927243e-15 pua1 = -1.104142481e-20
+ ub1 = -3.748327798e-19 lub1 = -8.960004008e-24 wub1 = -3.545141521e-25 pub1 = 5.630591775e-30
+ uc1 = 2.169604830e-10 luc1 = -2.166522453e-15 wuc1 = -1.564087500e-16 puc1 = 1.400177339e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.84 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 3.170859599e-01 lvth0 = 8.817240990e-07 wvth0 = 1.222905854e-07 pvth0 = -4.885553449e-13
+ k1 = -2.709787118e-01 lk1 = 1.221790345e-06 wk1 = 4.498077842e-07 pk1 = -6.467953404e-13
+ k2 = 4.031671796e-01 lk2 = -7.574489557e-07 wk2 = -2.430005125e-07 pk2 = 4.125360891e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.256182131e+00 ldsub = 7.284317864e-06 wdsub = 1.147703606e-06 pdsub = -4.603193557e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 2.240673878e-01 lvoff = -1.024825043e-06 wvoff = -1.959827088e-07 pvoff = 5.970682679e-13
+ nfactor = 1.364038402e+01 lnfactor = -3.413639107e-05 wnfactor = -6.376575489e-06 pnfactor = 1.996274622e-11
+ eta0 = -4.012882647e-01 leta0 = 1.930344234e-06 weta0 = 3.041414557e-07 peta0 = -1.219846292e-12
+ etab = 3.507488603e-01 letab = -1.687533639e-06 wetab = -2.658846688e-07 petab = 1.066406507e-12
+ u0 = 2.806354577e-02 lu0 = -1.338801750e-08 wu0 = 8.038198033e-10 pu0 = 3.286680199e-15
+ ua = 2.557894949e-09 lua = -1.639540283e-14 wua = -1.769021654e-15 pua = 9.201853888e-21
+ ub = -4.302580468e-18 lub = 2.595039055e-23 wub = 3.135343290e-24 pub = -1.508512560e-29
+ uc = -2.379563201e-10 luc = 6.272551334e-16 wuc = 1.481636926e-16 puc = -3.232055636e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 9.028145105e-01 la0 = 1.523651952e-06 wa0 = 3.871902937e-07 pa0 = -1.667491522e-12
+ ags = -1.000395022e+00 lags = 3.874668198e-06 wags = 7.185362784e-07 pags = -1.935297651e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.042275371e-07 lb0 = -3.819167856e-13 wb0 = -1.922511160e-13 pb0 = 2.413454382e-19
+ b1 = 4.089175861e-08 lb1 = -2.683227047e-13 wb1 = -2.584081080e-14 pb1 = 1.695617035e-19
+ keta = 1.969736027e-01 lketa = -5.817097006e-07 wketa = -1.064868830e-07 pketa = 3.201961399e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.179382640e+00 lpclm = 8.136197346e-06 wpclm = 2.330870809e-06 ppclm = -5.080544728e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -4.948768676e-03 lpdiblc2 = -2.199176451e-09 wpdiblc2 = 4.000513243e-09 ppdiblc2 = 6.364541126e-15
+ pdiblcb = 5.067425545e-02 lpdiblcb = -3.035132443e-07 wpdiblcb = -4.782098360e-08 ppdiblcb = 1.917997315e-13
+ drout = 0.56
+ pscbe1 = 1.101033985e+09 lpscbe1 = -6.053149235e+02 wpscbe1 = -2.596433974e+02 ppscbe1 = 5.220873084e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.227282992e-01 lkt1 = 9.748147854e-07 wkt1 = 1.434342517e-07 pkt1 = -6.108437850e-13
+ kt2 = -7.938462818e-02 lkt2 = 4.941245733e-07 wkt2 = 3.517995610e-08 pkt2 = -3.046095209e-13
+ at = 1.578766074e+05 lat = -7.169924669e-02 wat = 7.000991999e-03 pat = -2.807948069e-8
+ ute = -7.087306456e+00 lute = 2.923782047e-05 wute = 3.371484071e-06 pute = -1.678677282e-11
+ ua1 = -1.800301168e-08 lua1 = 8.907481063e-14 wua1 = 1.092717142e-14 pua1 = -5.079731497e-20
+ ub1 = 1.499778034e-17 lub1 = -7.061626550e-23 wub1 = -8.940876022e-24 pub1 = 4.006865175e-29
+ uc1 = -9.229235894e-11 luc1 = -9.261754840e-16 wuc1 = 5.435028445e-17 puc1 = 5.548679539e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.85 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 7.937800972e-01 lvth0 = -7.680579848e-08 wvth0 = -1.640195908e-07 pvth0 = 8.715314912e-14
+ k1 = 6.484758779e-01 lk1 = -6.270360717e-07 wk1 = -3.049074960e-08 pk1 = 3.189822272e-13
+ k2 = -1.005150039e-01 lk2 = 2.553481272e-07 wk2 = 3.104208571e-08 pk2 = -1.385049307e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.495600062e+00 ldsub = -4.281285244e-06 wdsub = -2.295407213e-06 pdsub = 2.320165475e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -3.198180790e-01 lvoff = 6.881223899e-08 wvoff = 1.388585976e-07 pvoff = -7.622594312e-14
+ nfactor = -6.058513806e+00 lnfactor = 5.473876890e-06 wnfactor = 5.572404867e-06 pnfactor = -4.064096199e-12
+ eta0 = 1.120880502e+00 leta0 = -1.130411413e-06 weta0 = -6.082827191e-07 peta0 = 6.148434642e-13
+ etab = -8.969676719e-01 letab = 8.213572965e-07 wetab = 5.317693376e-07 petab = -5.375050017e-13
+ u0 = 1.602787924e-02 lu0 = 1.081313225e-08 wu0 = 7.487636141e-09 pu0 = -1.015304412e-14
+ ua = -8.248751638e-09 lua = 5.334450837e-15 wua = 4.632663562e-15 pua = -3.670565122e-21
+ ub = 1.230099358e-17 lub = -7.435843687e-24 wub = -6.825140103e-24 pub = 4.943274956e-30
+ uc = -1.083141739e-10 luc = 3.665725207e-16 wuc = 9.237901644e-17 puc = -2.110345177e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.981918887e+04 lvsat = 1.009028725e-01 wvsat = 2.532338016e-02 pvsat = -5.091989829e-8
+ a0 = 7.116585410e+00 la0 = -1.097091158e-05 wa0 = -3.593451700e-06 pa0 = 6.336727671e-12
+ ags = 4.409992822e+00 lags = -7.004463935e-06 wags = -2.555445842e-06 pags = 4.647979762e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.401602900e-07 lb0 = -4.541698620e-13 wb0 = -2.149581724e-13 pb0 = 2.870044692e-19
+ b1 = 7.060957997e-10 lb1 = -1.875179366e-13 wb1 = -4.462045309e-16 pb1 = 1.184985847e-19
+ keta = -6.348267072e-01 lketa = 1.090862717e-06 wketa = 3.838371632e-07 pketa = -6.657405877e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.155315110e+00 lpclm = -2.590738205e-06 wpclm = -1.093786105e-06 ppclm = 1.805707450e-12
+ pdiblc1 = 5.371846616e-01 lpdiblc1 = -2.959568570e-07 wpdiblc1 = -6.024587525e-08 ppdiblc1 = 1.211415625e-13
+ pdiblc2 = -2.478774381e-02 lpdiblc2 = 3.769275700e-08 wpdiblc2 = 1.868584952e-08 ppdiblc2 = -2.316452746e-14
+ pdiblcb = 1.476230808e-01 lpdiblcb = -4.984565851e-07 wpdiblcb = -9.351813708e-08 ppdiblcb = 2.836869280e-13
+ drout = 3.904020436e+00 ldrout = -6.724109477e-06 wdrout = -2.009269098e-06 pdrout = 4.040210173e-12
+ pscbe1 = 3.976706747e+08 lpscbe1 = 8.089981747e+02 wpscbe1 = 2.542447752e+02 ppscbe1 = -5.112318345e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.345293063e-05 lalpha0 = -6.720636099e-11 walpha0 = -2.112025290e-11 palpha0 = 4.246830885e-17
+ alpha1 = 1.935871632e+00 lalpha1 = -2.183455474e-06 walpha1 = -5.884685850e-07 palpha1 = 1.183284392e-12
+ beta0 = 3.579543680e+01 lbeta0 = -4.410746922e-05 wbeta0 = -1.386170445e-05 pbeta0 = 2.787292124e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 7.346911206e-02 lkt1 = -2.240106225e-07 wkt1 = -2.531311393e-07 pkt1 = 1.865643512e-13
+ kt2 = 4.265088998e-01 lkt2 = -5.231190502e-07 wkt2 = -2.688742999e-07 pkt2 = 3.067785203e-13
+ at = 1.896562588e+04 lat = 2.076210102e-01 wat = 7.456434576e-02 pat = -1.639349266e-7
+ ute = 1.587559330e+01 lute = -1.693565688e-05 wute = -9.900478187e-06 pute = 9.900303079e-12
+ ua1 = 5.182949306e-08 lua1 = -5.134341226e-14 wua1 = -2.896074252e-14 pua1 = 2.940874395e-20
+ ub1 = -3.909037288e-17 lub1 = 3.814343576e-23 wub1 = 2.171600247e-23 pub1 = -2.157577033e-29
+ uc1 = -9.901999276e-10 luc1 = 8.793244844e-16 wuc1 = 5.758124179e-16 puc1 = -4.936808036e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.86 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 8.424746912e-01 lvth0 = -1.260256124e-07 wvth0 = -1.572711140e-07 pvth0 = 8.033188323e-14
+ k1 = -4.283618718e-01 lk1 = 4.614164500e-07 wk1 = 5.763252088e-07 pk1 = -2.943788481e-13
+ k2 = 3.152370518e-01 lk2 = -1.648882301e-07 wk2 = -2.142560502e-07 pk2 = 1.094389909e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -3.621758405e-01 lvoff = 1.116268713e-07 wvoff = 1.282607666e-07 pvoff = -6.551380394e-14
+ nfactor = -4.171259751e+00 lnfactor = 3.566266913e-06 wnfactor = 3.136825254e-06 pnfactor = -1.602246424e-12
+ eta0 = -4.954524662e-01 leta0 = 5.033553234e-07 weta0 = -3.846199902e-13 peta0 = 1.964585063e-19
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 3.501386970e-02 lu0 = -8.377641105e-09 wu0 = -5.169292668e-09 pu0 = 2.640402325e-15
+ ua = -4.378955446e-09 lua = 1.422915023e-15 wua = 2.024132699e-15 pua = -1.033898645e-21
+ ub = 8.328205928e-18 lub = -3.420205550e-24 wub = -3.910962216e-24 pub = 1.997664746e-30
+ uc = 4.605098122e-10 luc = -2.083868008e-16 wuc = -2.353182024e-16 puc = 1.201972433e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.317214727e+05 lvsat = 2.641859117e-01 wvsat = -5.064676031e-02 pvsat = 2.586965611e-8
+ a0 = -8.969601952e+00 la0 = 5.288781398e-06 wa0 = 5.409034001e-06 pa0 = -2.762858841e-12
+ ags = -5.253430486e+00 lags = 2.763189057e-06 wags = 4.129941761e-06 pags = -2.109516432e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.206812063e-07 lb0 = 1.127208706e-13 wb0 = 1.394555161e-13 pb0 = -7.123192522e-20
+ b1 = -3.736084496e-07 lb1 = 1.908339655e-13 wb1 = 2.360951348e-13 pb1 = -1.205940895e-19
+ keta = 9.056443002e-01 lketa = -4.662238103e-07 wketa = -5.555267136e-07 pketa = 2.837552680e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.285908178e+00 lpclm = 8.876021169e-07 wpclm = 1.400247536e-06 ppclm = -7.152268381e-13
+ pdiblc1 = 4.602994019e-01 lpdiblc1 = -2.182423128e-07 wpdiblc1 = 1.204917505e-07 ppdiblc1 = -6.154549928e-14
+ pdiblc2 = 2.522786576e-02 lpdiblc2 = -1.286232093e-08 wpdiblc2 = -8.554264740e-09 ppdiblc2 = 4.369398669e-15
+ pdiblcb = -6.018364499e-01 lpdiblcb = 2.590866161e-07 wpdiblcb = 3.783202085e-07 ppdiblcb = -1.932406660e-13
+ drout = -6.577532450e+00 ldrout = 3.870497439e-06 wdrout = 4.018538197e-06 pdrout = -2.052613051e-12
+ pscbe1 = 1.975543419e+09 lpscbe1 = -7.858935053e+02 wpscbe1 = -5.084895504e+02 ppscbe1 = 2.597293435e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.076934490e-05 lalpha0 = 3.814005601e-11 walpha0 = 4.224050580e-11 palpha0 = -2.157585900e-17
+ alpha1 = -1.321743263e+00 lalpha1 = 1.109296054e-06 walpha1 = 1.176937170e-06 palpha1 = -6.011630293e-13
+ beta0 = -3.425856997e+01 lbeta0 = 2.670214007e-05 wbeta0 = 2.772340889e-05 pbeta0 = -1.416072914e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.453106478e-02 lkt1 = -1.350612757e-07 wkt1 = -1.385941211e-07 pkt1 = 7.079193675e-14
+ kt2 = -1.465089572e-01 lkt2 = 5.607937740e-08 wkt2 = 7.000828446e-08 pkt2 = -3.575925159e-14
+ at = 4.426972833e+05 lat = -2.206810169e-01 wat = -1.771326595e-01 pat = 9.047688263e-8
+ ute = -4.391146268e-01 lute = -4.449785145e-07 wute = -2.139233308e-07 pute = 1.092690425e-13
+ ua1 = 1.240617085e-09 lua1 = -2.088846656e-16 wua1 = 2.712617097e-16 pua1 = -1.385566837e-22
+ ub1 = -2.091621868e-18 lub1 = 7.456162207e-25 wub1 = 7.489218910e-25 pub1 = -3.825388170e-31
+ uc1 = -2.489757399e-10 luc1 = 1.301054526e-16 wuc1 = 1.766846542e-16 puc1 = -9.024804776e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.87 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.375477052e-01 lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = 6.938893904e-24 pk2 = 8.673617380e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 7.806255642e-24 petab = 6.288372600e-30
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16
+ ub = 2.286030910e-18 lub = -3.339471417e-25 wub = -1.540743956e-39
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-07 wags = 2.220446049e-22 pags = -1.110223025e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = 1.387778781e-23 pketa = -3.469446952e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-07 wpclm = 4.440892099e-22
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = 1.387778781e-29
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 1.084202172e-25 ppdiblc2 = 5.692061406e-31
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-03 pat = 3.637978807e-24
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 wub1 = -7.703719778e-40
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = 4.523643975e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.88 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610889862e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456657017e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149736110e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935927057e-16
+ ags = 1.250000000e+00 lags = 6.286171583e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026246086e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347658096e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990252573e-18
+ drout = 5.033266586e-01 ldrout = 2.662110532e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629947662e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595196197e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865455e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275664625e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190826499e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.89 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 1.140963279e+00 lvth0 = -1.071407151e-07 wvth0 = -2.817473370e-07 pvth0 = 5.375344743e-14
+ k1 = 0.90707349
+ k2 = -1.379104027e-02 lk2 = -2.492342843e-08 wk2 = -5.259206361e-08 pk2 = 1.003382945e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999998e-03 lcdscd = 4.335403564e-19 wcdscd = 2.080779993e-18 pcdscd = -3.969845286e-25
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724287462e-17
+ nfactor = -1.367122711e+00 lnfactor = 6.277113832e-07 wnfactor = 1.783028553e-06 pnfactor = -3.401768854e-13
+ eta0 = 1.642889168e-09 leta0 = -2.641230358e-16 weta0 = 5.415415969e-19 peta0 = -1.033185551e-25
+ etab = -0.043998
+ u0 = -1.317993572e-01 lu0 = 3.008787420e-08 wu0 = 9.337280374e-08 pu0 = -1.781422373e-14
+ ua = 5.036359176e-10 lua = -3.045641810e-16 wua = -8.651215275e-16 pua = 1.650530758e-22
+ ub = -1.054947243e-17 lub = 2.284301680e-24 wub = 6.488611209e-24 pub = -1.237936178e-30
+ uc = 7.700399983e-11 luc = 2.675329576e-26 wuc = -1.431022460e-28 puc = 2.724526143e-35
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.500760136e+06 lvsat = -4.218004844e-01 wvsat = -1.254002619e+00 pvsat = 2.392461438e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.409772263e-06 lb0 = -8.442842676e-13 wb0 = -2.398208787e-12 pb0 = 4.575446617e-19
+ b1 = -3.020423958e-06 lb1 = 5.782830229e-13 wb1 = 1.642626163e-12 pb1 = -3.133900752e-19
+ keta = -2.700000009e-02 lketa = 1.436820107e-17 wketa = 8.160139231e-20 pketa = -1.557087792e-26
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.236013226e+00 lpclm = -2.016130945e-07 wpclm = -5.726866092e-07 ppclm = 1.092605874e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.200778689e-24 walpha0 = -1.631597215e-25 palpha0 = 3.112846081e-32
+ alpha1 = 0.85
+ beta0 = 1.005373824e+01 lbeta0 = 7.267793524e-07 wbeta0 = 2.064433393e-06 pbeta0 = -3.938649894e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.839584507e-02 lkt1 = -3.686397382e-08 wkt1 = -1.047129613e-07 pkt1 = 1.997776703e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.577747753e-11 wat = -3.469176590e-14 pat = 6.635673344e-21
+ ute = -2.268108645e+00 lute = 1.816948390e-07 wute = 5.161083492e-07 pute = -9.846624750e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.90 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.91 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = -1.525878906e-17
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-08 wkt1 = -1.776356839e-21
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.92 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-08 wketa = -5.551115123e-23 pketa = -2.220446049e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = -4.440892099e-22 ppclm = -3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267872e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.93 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15 wua1 = -6.617444900e-30 pua1 = -1.323488980e-35
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.94 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 weta0 = 3.469446952e-24 peta0 = 3.469446952e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -1.561251128e-22 petab = -2.949029909e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = 1.665334537e-22 pketa = -5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 5.929230631e-27 palpha0 = 1.312901068e-32
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.654361225e-30 pua1 = 4.963083675e-36
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = -1.540743956e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.95 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.522701748e-01 lvth0 = 2.220679177e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610700e-8
+ k2 = -8.011891576e-02 lk2 = 3.705406310e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026663e-01 lvoff = -9.262472634e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217668e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -2.498001805e-22 peta0 = -6.938893904e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.547523263e-02 lu0 = -3.505438827e-9
+ ua = -6.439246683e-10 lua = -4.848864078e-16
+ ub = 1.111503064e-18 lub = 2.659852385e-25
+ uc = 2.628890916e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.251774050e+05 lvsat = 3.119218935e-1
+ a0 = 1.011417809e+00 la0 = 1.906162389e-7
+ ags = 2.367344374e+00 lags = -1.129396050e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608784e-08 lb1 = -3.169227303e-14
+ keta = -1.194413445e-01 lketa = 5.737558588e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701757e-07 wpclm = 7.105427358e-21
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109111e-03 lpdiblc2 = -4.799688221e-9
+ pdiblcb = 9.625889888e-02 lpdiblcb = -9.749071472e-08 wpdiblcb = -1.422473250e-22 ppdiblcb = 1.066854938e-28
+ drout = 8.376749865e-01 ldrout = 8.291329324e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279453e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552323e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457427e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380072e-9
+ at = 1.158432509e+05 lat = -5.372855309e-2
+ ute = -8.338566439e-01 lute = -2.433498185e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563802e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648484e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475370e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.96 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.375477052e-01 lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = -2.220446049e-22 pk2 = 5.551115123e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-09 wcdscd = 5.551115123e-23
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 1.387778781e-23 petab = -5.204170428e-29
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16 wua = 1.323488980e-29
+ ub = 2.286030910e-18 lub = -3.339471417e-25
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-07 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = -5.551115123e-23 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-7
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = 2.220446049e-22 ppdiblc1 = -4.440892099e-28
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 2.125036258e-23 ppdiblc2 = 2.385244779e-30
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-03 pat = 2.910383046e-23
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 pub1 = 1.540743956e-45
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = -5.169878828e-32 puc1 = 1.421716678e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.97 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456612608e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149569577e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.936033638e-16
+ ags = 1.250000000e+00 lags = 6.285461041e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026379313e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990141551e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009866231e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.98 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = -3.567178047e+00 lvth0 = 7.911067358e-07 wvth0 = 2.269745108e-06 pvth0 = -4.330355901e-13
+ k1 = 0.90707349
+ k2 = -1.802308111e+00 lk2 = 3.163005895e-07 wk2 = 9.166625698e-07 pk2 = -1.748863850e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000027e-03 lcdscd = -5.141442827e-18 wcdscd = -1.375510816e-17 pcdscd = 2.624282736e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724220849e-17
+ nfactor = -1.367121211e+00 lnfactor = 6.277110970e-07 wnfactor = 1.783027739e-06 pnfactor = -3.401767303e-13
+ eta0 = 1.642889326e-09 leta0 = -2.641230346e-16 weta0 = 5.415449217e-19 peta0 = -1.033191894e-25
+ etab = -0.043998
+ u0 = 1.025634817e+00 lu0 = -1.907343621e-07 wu0 = -5.338778131e-07 pu0 = 1.018564124e-13
+ ua = 5.036486647e-10 lua = -3.045666130e-16 wua = -8.651284356e-16 pua = 1.650543937e-22
+ ub = -1.054935338e-17 lub = 2.284278967e-24 wub = 6.488546693e-24 pub = -1.237923869e-30
+ uc = 7.700399983e-11 luc = 2.713483281e-26 wuc = 9.429858983e-28 puc = -1.799117832e-34
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.989946961e+07 lvsat = 3.851849748e+00 wvsat = 1.088539869e+01 pvsat = -2.076781674e-6
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.409769924e-06 lb0 = -8.442838214e-13 wb0 = -2.398207520e-12 pb0 = 4.575444199e-19
+ b1 = -3.020424216e-06 lb1 = 5.782830722e-13 wb1 = 1.642626303e-12 pb1 = -3.133901019e-19
+ keta = -2.700000009e-02 lketa = 1.414912632e-17 wketa = -5.409006576e-19 pketa = 1.032507413e-25
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.236013822e+00 lpclm = -2.016132082e-07 wpclm = -5.726869319e-07 ppclm = 1.092606490e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.762597957e-24 walpha0 = 1.081661074e-24 palpha0 = -2.063584018e-31
+ alpha1 = 0.85
+ beta0 = 1.011879351e+01 lbeta0 = 7.143677172e-07 wbeta0 = 2.029177860e-06 pbeta0 = -3.871387271e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.440041678e-02 lkt1 = -3.571838560e-08 wkt1 = -1.014588917e-07 pkt1 = 1.935693611e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.587113366e-11 wat = 2.309679985e-13 pat = -4.423782229e-20
+ ute = -2.251844814e+00 lute = 1.785919276e-07 wute = 5.072944585e-07 pute = -9.678468056e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.99 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.100 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14 wb1 = 2.646977960e-29
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = -3.814697266e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.101 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647567e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 4.440892099e-22 ppclm = 2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267872e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.102 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-06 wpclm = 1.776356839e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.103 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159062e-03 leta0 = 4.128463499e-09 peta0 = -3.469446952e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = 1.734723476e-24 petab = -4.510281038e-29
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17 wuc = 1.033975766e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 pb0 = -5.293955920e-35
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = 1.387778781e-23 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = -7.411538288e-28 palpha0 = -1.799945013e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-02 wat = 2.328306437e-16
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -8.271806126e-31
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = 7.703719778e-46
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.104 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.522701748e-01 lvth0 = 2.220679177e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610700e-8
+ k2 = -8.011891576e-02 lk2 = 3.705406310e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026663e-01 lvoff = -9.262472634e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217668e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -4.024558464e-22 peta0 = -2.775557562e-29
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.547523263e-02 lu0 = -3.505438827e-9
+ ua = -6.439246683e-10 lua = -4.848864078e-16
+ ub = 1.111503064e-18 lub = 2.659852385e-25
+ uc = 2.628890916e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.251774050e+05 lvsat = 3.119218935e-1
+ a0 = 1.011417809e+00 la0 = 1.906162389e-7
+ ags = 2.367344374e+00 lags = -1.129396050e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608784e-08 lb1 = -3.169227303e-14
+ keta = -1.194413445e-01 lketa = 5.737558588e-08 pketa = -1.110223025e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701757e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109111e-03 lpdiblc2 = -4.799688221e-9
+ pdiblcb = 9.625889888e-02 lpdiblcb = -9.749071472e-08 wpdiblcb = -4.640385298e-23 ppdiblcb = 5.247538515e-29
+ drout = 8.376749865e-01 ldrout = 8.291329324e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279453e+02 wpscbe1 = 1.907348633e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552323e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457427e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380072e-9
+ at = 1.158432509e+05 lat = -5.372855309e-2
+ ute = -8.338566439e-01 lute = -2.433498185e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563802e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648484e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475370e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.105 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.375477052e-01 lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = -8.326672685e-23 pk2 = 3.469446952e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 1.561251128e-23 petab = 9.540979118e-30
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16
+ ub = 2.286030910e-18 lub = -3.339471417e-25
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = -2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-7
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = -8.326672685e-29
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = -1.951563910e-24 ppdiblc2 = 1.219727444e-30
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-03 pat = 7.275957614e-24
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 wub1 = -1.540743956e-39 pub1 = -3.851859889e-46
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = -3.877409121e-32 puc1 = -6.462348536e-39
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.106 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610978680e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456701426e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149680599e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.286171583e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026290495e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347671974e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990141551e-18
+ drout = 5.033266586e-01 ldrout = 2.662110532e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009864680e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190826499e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.107 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 1.625879187e+00 lvth0 = -1.996558816e-07 wvth0 = -4.926082127e-07 pvth0 = 9.398275046e-14
+ k1 = 0.90707349
+ k2 = 2.979877433e-01 lk2 = -8.440645544e-08 wk2 = -2.005520048e-07 pk2 = 3.826251479e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584979911e-01 ldsub = 2.518544814e-11 wdsub = 7.021975303e-11 pdsub = -1.339694580e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079655892e-19
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724309667e-17
+ nfactor = 1.334758346e+01 lnfactor = -2.179648549e-06 wnfactor = -6.044194547e-06 pnfactor = 1.153147701e-12
+ eta0 = 1.826783307e-02 leta0 = -3.485246401e-09 weta0 = -9.717243132e-09 peta0 = 1.853913948e-15
+ etab = -0.043998
+ u0 = -3.317912352e-01 lu0 = 6.824352463e-08 wu0 = 1.881805416e-07 pu0 = -3.590221282e-14
+ ua = -3.087980150e-09 lua = 3.806658820e-16 wua = 1.045373863e-15 pua = -1.994426978e-22
+ ub = 2.653989546e-17 lub = -4.791830462e-24 wub = -1.324041162e-23 pub = 2.526085172e-30
+ uc = 3.575979994e-10 luc = -5.353340678e-17 wuc = -1.492569274e-16 puc = 2.847613215e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.124878107e+07 lvsat = -2.090800406e+00 wvsat = -5.683352593e+00 pvsat = 1.084304108e-6
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325206324e-05 lb0 = 2.525346681e-12 wb0 = 6.996686721e-12 pb0 = -1.334869873e-18
+ b1 = 2.663302983e-06 lb1 = -5.060925053e-13 wb1 = -1.380730074e-12 pb1 = 2.634239678e-19
+ keta = -2.700000009e-02 lketa = 1.434302677e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564203824e-01 lpclm = 1.022009439e-07 wpclm = 2.743797791e-07 ppclm = -5.234782053e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150539047e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091395e-01 lkt1 = 5.088104398e-08 wkt1 = 1.399896830e-07 pkt1 = -2.670807166e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578824595e-11
+ ute = 4.121252916e-01 lute = -3.296562729e-07 wute = -9.097564876e-07 pute = 1.735688012e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.108 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.109 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.110 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 1.332267630e-21
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.111 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-01 wat = -9.313225746e-16
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.112 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159062e-03 leta0 = 4.128463499e-09 peta0 = -6.938893904e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -1.873501354e-22 petab = 1.734723476e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15 pua = -3.308722450e-36
+ ub = -2.930959084e-19 lub = 1.685734216e-24 pub = -3.081487911e-45
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -2.775557562e-23 pketa = 2.220446049e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 7.623296525e-27 palpha0 = -6.988021815e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.654361225e-30
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = 1.540743956e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.113 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.522701748e-01 lvth0 = 2.220679177e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610700e-8
+ k2 = -8.011891576e-02 lk2 = 3.705406310e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026663e-01 lvoff = -9.262472634e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217668e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 4.718447855e-22 peta0 = 6.245004514e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.547523263e-02 lu0 = -3.505438827e-9
+ ua = -6.439246683e-10 lua = -4.848864078e-16
+ ub = 1.111503064e-18 lub = 2.659852385e-25
+ uc = 2.628890916e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.251774050e+05 lvsat = 3.119218935e-01 wvsat = 4.656612873e-16 pvsat = -4.656612873e-22
+ a0 = 1.011417809e+00 la0 = 1.906162389e-7
+ ags = 2.367344374e+00 lags = -1.129396050e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608784e-08 lb1 = -3.169227303e-14
+ keta = -1.194413445e-01 lketa = 5.737558588e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701757e-07 wpclm = -7.105427358e-21
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109111e-03 lpdiblc2 = -4.799688221e-9
+ pdiblcb = 9.625889888e-02 lpdiblcb = -9.749071472e-08 wpdiblcb = -3.122502257e-23 ppdiblcb = 1.847480502e-28
+ drout = 8.376749865e-01 ldrout = 8.291329324e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279453e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552323e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457427e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380072e-9
+ at = 1.158432509e+05 lat = -5.372855309e-2
+ ute = -8.338566439e-01 lute = -2.433498185e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563802e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648484e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475370e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.114 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.375477052e-01 lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = 5.551115123e-23 pk2 = -8.326672685e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 2.775557562e-23 petab = -3.816391647e-29
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16
+ ub = 2.286030910e-18 lub = -3.339471417e-25
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-07 wags = 1.776356839e-21 pags = 8.881784197e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = -1.110223025e-22 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-7
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = 4.440892099e-22 ppdiblc1 = -5.551115123e-29
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 1.301042607e-23 ppdiblc2 = -1.084202172e-31
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-3
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 wub1 = 6.162975822e-39 pub1 = -1.540743956e-45
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = 2.067951531e-31 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.115 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456612608e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016978168e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149569577e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.286171583e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-08 wketa = -8.881784197e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026379313e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990585640e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.630233765e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865197e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.116 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 8.061145465e-01 lvth0 = -4.325626486e-08 wvth0 = -8.114210699e-08 pvth0 = 1.548077803e-14
+ k1 = 0.90707349
+ k2 = -1.872942668e-01 lk2 = 8.178558149e-09 wk2 = 4.302656511e-08 pk2 = -8.208866250e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584992040e-01 ldsub = 2.495405448e-11 wdsub = 6.961098779e-11 pdsub = -1.328080192e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079725281e-19
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724220849e-17
+ nfactor = 1.334758330e+01 lnfactor = -2.179648517e-06 wnfactor = -6.044194464e-06 pnfactor = 1.153147685e-12
+ eta0 = 1.826779867e-02 leta0 = -3.485240187e-09 weta0 = -9.717226783e-09 peta0 = 1.853910829e-15
+ etab = -0.043998
+ u0 = -8.465704720e-02 lu0 = 2.109378145e-08 wu0 = 6.413598440e-08 pu0 = -1.223624792e-14
+ ua = -3.087979294e-09 lua = 3.806657188e-16 wua = 1.045373434e-15 pua = -1.994426159e-22
+ ub = 2.653968253e-17 lub = -4.791789839e-24 wub = -1.324030475e-23 pub = 2.526064782e-30
+ uc = 3.550112941e-10 luc = -5.303989961e-17 wuc = -1.479585772e-16 puc = 2.822842511e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.914970573e+05 lvsat = 1.490802965e-01 wvsat = 2.094686876e-01 pvsat = -3.996369303e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325212843e-05 lb0 = 2.525359119e-12 wb0 = 6.996719441e-12 pb0 = -1.334876115e-18
+ b1 = 2.663317764e-06 lb1 = -5.060953252e-13 wb1 = -1.380737492e-12 pb1 = 2.634253832e-19
+ keta = -2.700000009e-02 lketa = 1.434297126e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564208446e-01 lpclm = 1.022010321e-07 wpclm = 2.743800111e-07 ppclm = -5.234786480e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150327289e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091288e-01 lkt1 = 5.088104192e-08 wkt1 = 1.399896776e-07 pkt1 = -2.670807063e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578778028e-11
+ ute = 3.963587508e-01 lute = -3.266482377e-07 wute = -9.018427563e-07 pute = 1.720589721e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.117 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.118 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = 7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.119 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-07 pk2 = 2.220446049e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647567e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 4.440892099e-22 ppclm = -2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15 wua1 = 3.308722450e-30
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16 wuc1 = -5.169878828e-32 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.120 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-06 wdsub = -1.776356839e-21
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14 wb0 = -1.058791184e-28
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14 pb1 = 2.646977960e-35
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.121 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 weta0 = -1.734723476e-24
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -3.295974604e-23 petab = 4.163336342e-29
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24 pub = -1.540743956e-45
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-06 pags = -1.776356839e-27
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = 5.293955920e-29 pb0 = 5.293955920e-35
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = 2.775557562e-23 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 7.411538288e-28 palpha0 = 4.976318565e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.240770919e-30 pua1 = -8.271806126e-37
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = -7.703719778e-46
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.122 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.821975320e-01 lvth0 = 9.303523806e-08 wvth0 = 3.447097530e-08 pvth0 = -3.484277924e-14
+ k1 = 6.351021960e-01 lk1 = -8.178610772e-08 wk1 = -3.526778869e-16 pk1 = 3.564819551e-22
+ k2 = -9.819090370e-02 lk2 = 5.532097549e-08 wk2 = 8.890189169e-09 pk2 = -8.986078750e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076448e-01 ldsub = 5.194667313e-08 wdsub = -1.040207920e-16 pdsub = 1.051430054e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026654e-01 lvoff = -9.262473516e-09 wvoff = -4.291291766e-16 pvoff = 4.337576964e-22
+ nfactor = 1.616966924e+00 lnfactor = 6.097217582e-07 wnfactor = -4.169514511e-15 pnfactor = 4.214484761e-21
+ eta0 = -4.954531764e-01 leta0 = 5.033556864e-07 weta0 = 2.379968514e-16 peta0 = -2.405640999e-22
+ etab = -1.699316551e-01 letab = 8.647946918e-08 wetab = 4.781841589e-17 petab = -4.833422551e-23
+ u0 = -2.210078630e-03 lu0 = 2.447848620e-08 wu0 = 1.361929054e-08 pu0 = -1.376618821e-14
+ ua = -6.439294864e-10 lua = -4.848815377e-16 wua = 2.370166855e-21 pua = -2.395731474e-27
+ ub = 1.111498246e-18 lub = 2.659901090e-25 wub = 2.370352916e-30 pub = -2.395919541e-36
+ uc = 2.628890927e-11 luc = 1.340715722e-17 wuc = -5.360678376e-26 puc = 5.418487962e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.914931349e+06 lvsat = 3.030687524e+00 wvsat = 1.323176037e+00 pvsat = -1.337447814e-6
+ a0 = 1.011417803e+00 la0 = 1.906162443e-07 wa0 = 2.592706494e-15 pa0 = -2.620669903e-21
+ ags = 2.367344351e+00 lags = -1.129396027e-06 wags = 1.145646067e-14 pags = -1.158003116e-20
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907885e-08 lb0 = -1.871983642e-14 wb0 = -2.718684593e-23 pb0 = 2.748010462e-29
+ b1 = 6.204608816e-08 lb1 = -3.169227335e-14 wb1 = -1.572521961e-22 pb1 = 1.589483266e-28
+ keta = -1.194413453e-01 lketa = 5.737558669e-08 wketa = 3.952973504e-16 pketa = -3.995610509e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898536e+00 lpclm = -4.321701819e-07 wpclm = -3.028485906e-15 ppclm = 3.061151332e-21
+ pdiblc1 = 6.826367982e-01 lpdiblc1 = -3.318091416e-07 wpdiblc1 = 5.676632497e-16 ppdiblc1 = -5.737854636e-22
+ pdiblc2 = 9.443109138e-03 lpdiblc2 = -4.799688249e-09 wpdiblc2 = -1.368019587e-17 ppdiblc2 = 1.382775838e-23
+ pdiblcb = 9.625889866e-02 lpdiblcb = -9.749071449e-08 wpdiblcb = 1.099100186e-16 ppdiblcb = -1.110955247e-22
+ drout = 8.376749873e-01 ldrout = 8.291329245e-08 wdrout = -3.815046057e-16 pdrout = 3.856222008e-22
+ pscbe1 = 1.037253089e+09 lpscbe1 = -3.066279363e+02 wpscbe1 = 4.392906189e-06 ppscbe1 = -4.440286636e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946629e-06 lalpha0 = -1.672796883e-12 walpha0 = 5.156357112e-21 palpha0 = -5.211976684e-27
+ alpha1 = 0.85
+ beta0 = 1.689804916e+01 lbeta0 = 5.720551851e-07 wbeta0 = -2.295894319e-14 pbeta0 = 2.320655312e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718610e-01 lkt1 = -4.432457352e-09 wkt1 = 3.684341721e-17 pkt1 = -3.724087705e-23
+ kt2 = -1.732617330e-02 lkt2 = -9.905380060e-09 wkt2 = 6.005085318e-18 pkt2 = -6.069811320e-24
+ at = 1.158432499e+05 lat = -5.372855215e-02 wat = 4.562644754e-10 pat = -4.611859331e-16
+ ute = -8.338566420e-01 lute = -2.433498205e-07 wute = -9.430962677e-16 pute = 9.532676870e-22
+ ua1 = 1.741162740e-09 lua1 = -4.645563762e-16 wua1 = 1.953780755e-24 pua1 = -1.974854008e-30
+ ub1 = -7.096737815e-19 lub1 = 3.973648573e-26 wub1 = 4.286565388e-34 pub1 = -4.332787707e-40
+ uc1 = 7.705161076e-11 luc1 = -3.642475380e-17 wuc1 = -4.747582446e-26 puc1 = 4.798784926e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.123 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 7.776929907e-01 lvth0 = -5.789970531e-08 wvth0 = -6.894195061e-08 pvth0 = 1.797909553e-14
+ k1 = 2.425254185e-02 lk1 = 2.302273437e-07 wk1 = 7.053557738e-16 pk1 = -1.839470798e-22
+ k2 = 1.741672963e-01 lk2 = -8.379578003e-08 wk2 = -1.778037834e-08 pk2 = 4.636873745e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850176e-01 ldsub = 7.902988878e-08 wdsub = 2.080424721e-16 pdsub = -5.425460081e-23
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895709e-01 lvoff = -1.856546724e-08 wvoff = 8.582583533e-16 pvoff = -2.238217389e-22
+ nfactor = 4.181852111e+00 lnfactor = -7.003856872e-07 wnfactor = 8.339029023e-15 pnfactor = -2.174701308e-21
+ eta0 = 1.000416473e+00 leta0 = -2.607135883e-07 weta0 = -4.759943550e-16 peta0 = 1.241322600e-22
+ etab = 4.461928492e-02 letab = -2.311014727e-08 wetab = -9.563704863e-17 petab = 2.494078381e-23
+ u0 = 7.223690378e-02 lu0 = -1.354799016e-08 wu0 = -2.723858107e-08 pu0 = 7.103440604e-15
+ ua = -2.102021197e-09 lua = 2.598912947e-16 wua = -4.740333710e-21 pua = 1.236212667e-27
+ ub = 2.286040547e-18 lub = -3.339496549e-25 wub = -4.740705826e-30 pub = 1.236309710e-36
+ uc = 1.078724744e-11 luc = 2.132518905e-17 wuc = 1.072133607e-25 puc = -2.795979038e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.882720731e+06 lvsat = -1.463029992e+00 wvsat = -2.646352074e+00 pvsat = 6.901315721e-7
+ a0 = 1.264221194e+00 la0 = 6.148781164e-08 wa0 = -5.185412988e-15 pa0 = 1.352281842e-21
+ ags = -9.846887014e-01 lags = 5.827755276e-07 wags = -2.291292400e-14 pags = 5.975369533e-21
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.152151564e-16 lb0 = 3.004649978e-23 wb0 = 5.437371919e-23 pb0 = -1.417990473e-29
+ b1 = -6.664189737e-16 lb1 = 1.737927385e-22 wb1 = 3.145044391e-22 pb1 = -8.201835465e-29
+ keta = 7.220181600e-02 lketa = -4.051305711e-08 wketa = -7.905947008e-16 pketa = 2.061760276e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500137e-01 lpclm = -1.136192480e-07 wpclm = 6.056973589e-15 ppclm = -1.579573805e-21
+ pdiblc1 = -3.048846444e-01 lpdiblc1 = 1.726029860e-07 wpdiblc1 = -1.135325833e-15 ppdiblc1 = 2.960770240e-22
+ pdiblc2 = -8.673906618e-03 lpdiblc2 = 4.454229761e-09 wpdiblc2 = 2.736040409e-17 ppdiblc2 = -7.135207789e-24
+ pdiblcb = -8.553970401e-02 lpdiblcb = -4.630533427e-09 wpdiblcb = -2.198201621e-16 ppdiblcb = 5.732603281e-23
+ drout = 1.518101609e+00 ldrout = -2.646391000e-07 wdrout = 7.630127641e-16 pdrout = -1.989830523e-22
+ pscbe1 = 6.718078115e+07 lpscbe1 = 1.888714176e+02 wpscbe1 = -8.785812378e-06 ppscbe1 = 2.291216850e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729711e-06 lalpha0 = -2.066502091e-12 walpha0 = -1.031272778e-20 palpha0 = 2.689410923e-27
+ alpha1 = 0.85
+ beta0 = 2.187554641e+01 lbeta0 = -1.970380727e-06 wbeta0 = 4.591782954e-14 pbeta0 = -1.197473409e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774103e-01 lkt1 = 2.024134099e-08 wkt1 = -7.368683441e-17 pkt1 = 1.921640624e-23
+ kt2 = -4.489649531e-02 lkt2 = 4.177154438e-09 wkt2 = -1.201017064e-17 pkt2 = 3.132077930e-24
+ at = -8.189371221e+03 lat = 9.625574286e-03 wat = -9.125292418e-10 pat = 2.379748476e-16
+ ute = -1.301136477e+00 lute = -4.669822644e-09 wute = 1.886192535e-15 pute = -4.918909724e-22
+ ua1 = 1.724096906e-09 lua1 = -4.558393872e-16 wua1 = -3.907558200e-24 pua1 = 1.019036057e-30
+ ub1 = -2.029308258e-18 lub1 = 7.137873014e-25 wub1 = -8.573099962e-34 pub1 = 2.235750443e-40
+ uc1 = -1.418079326e-10 luc1 = 7.536563689e-17 wuc1 = 9.495149383e-26 puc1 = -2.476198768e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.124 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456790244e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149680599e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935927057e-16
+ ags = 1.250000000e+00 lags = 6.285816312e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026201677e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347671974e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662101650e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.630043030e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865197e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.191033295e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.125 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 9.627035343e-01 lvth0 = -7.313125148e-08 wvth0 = -1.581732409e-07 pvth0 = 3.017723995e-14
+ k1 = 0.90707349
+ k2 = -4.976247873e-01 lk2 = 6.738527684e-08 wk2 = 1.956880787e-07 pk2 = -3.733454579e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585002188e-01 ldsub = 2.476043415e-11 wdsub = 6.911174762e-11 pdsub = -1.318555388e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079655892e-19
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724309667e-17
+ nfactor = 1.334758404e+01 lnfactor = -2.179648659e-06 wnfactor = -6.044194829e-06 pnfactor = 1.153147755e-12
+ eta0 = 1.826779849e-02 leta0 = -3.485240153e-09 weta0 = -9.717226695e-09 peta0 = 1.853910812e-15
+ etab = -0.043998
+ u0 = 4.637763925e-01 lu0 = -8.353964079e-08 wu0 = -2.056559745e-07 pu0 = 3.923628075e-14
+ ua = -3.087976251e-09 lua = 3.806651381e-16 wua = 1.045371936e-15 pua = -1.994423302e-22
+ ub = 2.653990193e-17 lub = -4.791831698e-24 wub = -1.324041268e-23 pub = 2.526085373e-30
+ uc = 3.528542115e-10 luc = -5.262835845e-17 wuc = -1.468974392e-16 puc = 2.802597484e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.016421737e+06 lvsat = 1.203158576e+00 wvsat = 2.927355935e+00 pvsat = -5.584985294e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325201989e-05 lb0 = 2.525338411e-12 wb0 = 6.996666048e-12 pb0 = -1.334865929e-18
+ b1 = 2.663305599e-06 lb1 = -5.060930044e-13 wb1 = -1.380731508e-12 pb1 = 2.634242415e-19
+ keta = -2.700000009e-02 lketa = 1.434308228e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564201645e-01 lpclm = 1.022009023e-07 wpclm = 2.743796765e-07 ppclm = -5.234780096e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150539047e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091390e-01 lkt1 = 5.088104389e-08 wkt1 = 1.399896827e-07 pkt1 = -2.670807160e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578824595e-11
+ ute = 3.832108188e-01 lute = -3.241397963e-07 wute = -8.953748678e-07 pute = 1.708249895e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.126 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.127 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-07 wa0 = 1.776356839e-21
+ ags = 3.207608585e-01 lags = 4.826429794e-07 wags = -4.440892099e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.128 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-07 pk2 = -1.110223025e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-08 pketa = -5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 ppclm = 3.108624469e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.129 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.130 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 weta0 = 8.673617380e-25
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -4.336808690e-24 petab = -6.938893904e-30
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15 pua = 8.271806126e-37
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-06 pags = 8.881784197e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = 5.293955920e-29 pb0 = 5.293955920e-35
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 2.805796638e-27 palpha0 = -1.799945013e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = 4.135903063e-31 pua1 = -1.654361225e-36
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 wub1 = -3.851859889e-40 pub1 = -3.851859889e-46
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.131 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.552397824e-01 lvth0 = 1.920515398e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610696e-8
+ k2 = -7.935304322e-02 lk2 = 3.627992986e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667335e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026664e-01 lvoff = -9.262472597e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217672e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -7.632783294e-23 peta0 = 1.214306433e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.664850807e-02 lu0 = -4.691369216e-9
+ ua = -6.439244642e-10 lua = -4.848866142e-16
+ ub = 1.111503269e-18 lub = 2.659850321e-25
+ uc = 2.628890915e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111883581e+05 lvsat = 1.967033607e-01 pvsat = 1.164153218e-22
+ a0 = 1.011417809e+00 la0 = 1.906162387e-7
+ ags = 2.367344375e+00 lags = -1.129396051e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608782e-08 lb1 = -3.169227302e-14
+ keta = -1.194413445e-01 lketa = 5.737558585e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701755e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109109e-03 lpdiblc2 = -4.799688220e-9
+ pdiblcb = 9.625889889e-02 lpdiblcb = -9.749071473e-08 wpdiblcb = -1.908195824e-23 ppdiblcb = -2.146720302e-29
+ drout = 8.376749865e-01 ldrout = 8.291329327e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279457e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552343e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457430e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380073e-9
+ at = 1.158432509e+05 lat = -5.372855313e-2
+ ute = -8.338566440e-01 lute = -2.433498184e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563804e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648481e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475369e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.132 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.316084900e-01 lvth0 = -1.980291269e-8
+ k1 = 2.425254334e-02 lk1 = 2.302273434e-7
+ k2 = 1.364915753e-01 lk2 = -7.397047947e-08 wk2 = 2.775557562e-23 pk2 = 5.204170428e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988866e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546771e-8
+ nfactor = 4.181852129e+00 lnfactor = -7.003856918e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928472e-02 letab = -2.311014721e-08 wetab = -6.938893904e-24 petab = 1.214306433e-29
+ u0 = 1.451973038e-02 lu0 = 1.503840623e-9
+ ua = -2.102031242e-09 lua = 2.598939142e-16
+ ub = 2.286030502e-18 lub = -3.339470352e-25
+ uc = 1.078724767e-11 luc = 2.132518899e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.752347497e+05 lvsat = -6.761528150e-4
+ a0 = 1.264221183e+00 la0 = 6.148781451e-8
+ ags = -9.846887499e-01 lags = 5.827755403e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.220181432e-02 lketa = -4.051305667e-08 wketa = 1.387778781e-23 pketa = -1.734723476e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500265e-01 lpclm = -1.136192514e-7
+ pdiblc1 = -3.048846468e-01 lpdiblc1 = 1.726029866e-07 ppdiblc1 = 6.938893904e-29
+ pdiblc2 = -8.673906560e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 3.252606517e-25 ppdiblc2 = -3.523657061e-31
+ pdiblcb = -8.553970447e-02 lpdiblcb = -4.630533306e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076254e+07 lpscbe1 = 1.888714225e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729689e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380753e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-08 wkt1 = 4.440892099e-22
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373154e+03 lat = 9.625574790e-3
+ ute = -1.301136473e+00 lute = -4.669823687e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393851e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873019e-25
+ uc1 = -1.418079323e-10 luc1 = 7.536563684e-17 wuc1 = 5.169878828e-32 puc1 = 2.261821987e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.133 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456701426e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149680599e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.285993948e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026201677e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347658096e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.630043030e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009864680e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190826499e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.134 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 1.640247921e+00 lvth0 = -2.023972348e-07 wvth0 = -4.779281183e-07 pvth0 = 9.118199398e-14
+ k1 = 0.90707349
+ k2 = -3.443785481e-01 lk2 = 3.814803985e-08 wk2 = 1.233662746e-07 pk2 = -2.353655806e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585021073e-01 ldsub = 2.440014616e-11 wdsub = 6.822053216e-11 pdsub = -1.301552245e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079517114e-19
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724309667e-17
+ nfactor = 1.334758347e+01 lnfactor = -2.179648551e-06 wnfactor = -6.044194562e-06 pnfactor = 1.153147704e-12
+ eta0 = 1.826777218e-02 leta0 = -3.485235134e-09 weta0 = -9.717214281e-09 peta0 = 1.853908444e-15
+ etab = -0.043998
+ u0 = 2.066270621e-01 lu0 = -3.447914862e-08 wu0 = -8.429897664e-08 pu0 = 1.608306456e-14
+ ua = -3.087977982e-09 lua = 3.806654685e-16 wua = 1.045372754e-15 pua = -1.994424862e-22
+ ub = 2.653983749e-17 lub = -4.791819404e-24 wub = -1.324038227e-23 pub = 2.526079571e-30
+ uc = 3.488330108e-10 luc = -5.186116966e-17 wuc = -1.449997060e-16 puc = 2.766391390e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.128720330e+06 lvsat = 8.430115758e-01 wvsat = 2.036489235e+00 pvsat = -3.885336351e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325205743e-05 lb0 = 2.525345573e-12 wb0 = 6.996683763e-12 pb0 = -1.334869308e-18
+ b1 = 2.663308614e-06 lb1 = -5.060935796e-13 wb1 = -1.380732931e-12 pb1 = 2.634245130e-19
+ keta = -2.700000009e-02 lketa = 1.434302677e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564203852e-01 lpclm = 1.022009444e-07 wpclm = 2.743797807e-07 ppclm = -5.234782084e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150539047e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091505e-01 lkt1 = 5.088104606e-08 wkt1 = 1.399896881e-07 pkt1 = -2.670807262e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578801312e-11
+ ute = 3.587006802e-01 lute = -3.194636050e-07 wute = -8.838077490e-07 pute = 1.686181452e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.135 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.136 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-07 wvth0 = 1.776356839e-21
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = 7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.137 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647567e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = -4.440892099e-22 ppclm = -7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-08 ppdiblc2 = -2.775557562e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267872e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.138 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14 wb0 = 2.117582368e-28
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-06 wpclm = -3.552713679e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.139 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 peta0 = 3.469446952e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -1.734723476e-23 petab = 1.075528555e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24 pub = -3.081487911e-45
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = -1.058791184e-28 pb0 = -1.058791184e-34
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -1.110223025e-22 pketa = -1.665334537e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 6.564505341e-27 palpha0 = -4.235164736e-34
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.654361225e-30
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 wub1 = -7.703719778e-40 pub1 = 2.311115933e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.140 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.552397824e-01 lvth0 = 1.920515398e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610696e-8
+ k2 = -7.935304322e-02 lk2 = 3.627992986e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667335e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026664e-01 lvoff = -9.262472597e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217672e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 2.498001805e-22 peta0 = -1.387778781e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.664850807e-02 lu0 = -4.691369216e-9
+ ua = -6.439244642e-10 lua = -4.848866142e-16
+ ub = 1.111503269e-18 lub = 2.659850321e-25
+ uc = 2.628890915e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111883581e+05 lvsat = 1.967033607e-1
+ a0 = 1.011417809e+00 la0 = 1.906162387e-7
+ ags = 2.367344375e+00 lags = -1.129396051e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608782e-08 lb1 = -3.169227302e-14
+ keta = -1.194413445e-01 lketa = 5.737558585e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701755e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109109e-03 lpdiblc2 = -4.799688220e-9
+ pdiblcb = 9.625889889e-02 lpdiblcb = -9.749071473e-08 wpdiblcb = 1.023486851e-22 ppdiblcb = 6.028164079e-29
+ drout = 8.376749865e-01 ldrout = 8.291329327e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279457e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552343e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457430e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380073e-9
+ at = 1.158432509e+05 lat = -5.372855313e-2
+ ute = -8.338566440e-01 lute = -2.433498184e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563804e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648481e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475369e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.141 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.316084900e-01 lvth0 = -1.980291269e-8
+ k1 = 2.425254334e-02 lk1 = 2.302273434e-7
+ k2 = 1.364915753e-01 lk2 = -7.397047947e-08 wk2 = -1.665334537e-22 pk2 = -9.714451465e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988866e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546771e-8
+ nfactor = 4.181852129e+00 lnfactor = -7.003856918e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928472e-02 letab = -2.311014721e-08 wetab = 4.857225733e-23 petab = -1.387778781e-29
+ u0 = 1.451973038e-02 lu0 = 1.503840623e-9
+ ua = -2.102031242e-09 lua = 2.598939142e-16
+ ub = 2.286030502e-18 lub = -3.339470352e-25
+ uc = 1.078724767e-11 luc = 2.132518899e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.752347497e+05 lvsat = -6.761528150e-4
+ a0 = 1.264221183e+00 la0 = 6.148781451e-8
+ ags = -9.846887499e-01 lags = 5.827755403e-07 wags = 1.776356839e-21 pags = -4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.220181432e-02 lketa = -4.051305667e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500265e-01 lpclm = -1.136192514e-7
+ pdiblc1 = -3.048846468e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = 4.440892099e-22 ppdiblc1 = -1.110223025e-28
+ pdiblc2 = -8.673906560e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = -4.119968255e-24 ppdiblc2 = -5.854691731e-30
+ pdiblcb = -8.553970447e-02 lpdiblcb = -4.630533306e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076254e+07 lpscbe1 = 1.888714225e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729689e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380753e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373154e+03 lat = 9.625574790e-03 pat = 1.455191523e-23
+ ute = -1.301136473e+00 lute = -4.669823687e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393851e-16 wua1 = -6.617444900e-30
+ ub1 = -2.029308260e-18 lub1 = 7.137873019e-25 pub1 = -7.703719778e-46
+ uc1 = -1.418079323e-10 luc1 = 7.536563684e-17 wuc1 = -2.584939414e-32 puc1 = 6.462348536e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.142 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456790244e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.150013666e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935820476e-16
+ ags = 1.250000000e+00 lags = 6.286882126e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026379313e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990585640e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009866231e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.143 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = -2.712151192e+00 lvth0 = 6.279795823e-07 wvth0 = 1.445536326e-06 pvth0 = -2.757880936e-13
+ k1 = 0.90707349
+ k2 = 2.080083157e-01 lk2 = -6.723964035e-08 wk2 = -1.207511569e-07 pk2 = 2.303763022e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.687830613e+00 ldsub = -4.253002681e-07 wdsub = -9.851433845e-07 pdsub = 1.879515657e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079586503e-19
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724220849e-17
+ nfactor = -3.997886150e+00 lnfactor = 1.129624217e-06 wnfactor = 1.621323520e-06 pnfactor = -3.093258290e-13
+ eta0 = -1.264688194e-02 leta0 = 2.412848068e-09 weta0 = 3.944960646e-09 peta0 = -7.526432618e-16
+ etab = -0.043998
+ u0 = 4.427431561e-01 lu0 = -7.952679374e-08 wu0 = -1.886462343e-07 pu0 = 3.599106046e-14
+ ua = -1.023251079e-09 lua = -1.325551842e-17 wua = 1.329038639e-16 pua = -2.535619658e-23
+ ub = -4.555577596e-18 lub = 1.140750460e-24 wub = 5.016767147e-25 pub = -9.571289368e-32
+ uc = -2.391896018e-10 luc = 6.032531251e-17 wuc = 1.148663033e-16 puc = -2.191488254e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.313909858e+06 lvsat = -9.585100672e-01 wvsat = -2.136511210e+00 pvsat = 4.076164276e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.404797633e-06 lb0 = -6.525491778e-13 wb0 = -3.645135095e-13 pb0 = 6.954407442e-20
+ b1 = 2.644971507e-06 lb1 = -5.025951163e-13 wb1 = -1.372629177e-12 pb1 = 2.618784301e-19
+ keta = -8.680480736e-01 lketa = 1.604601978e-07 wketa = 3.716860572e-07 pketa = -7.091249611e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.238634796e-02 lpclm = 3.183778305e-08 wpclm = 1.113922835e-07 ppclm = -2.125208819e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.999997308e-08 lalpha0 = 5.135634875e-21 walpha0 = 1.190335528e-20 palpha0 = -2.270993587e-27
+ alpha1 = 0.85
+ beta0 = 1.393352495e+01 lbeta0 = -1.342963468e-08 wbeta0 = 1.137225354e-13 pbeta0 = -2.169667823e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.815416568e-01 lkt1 = -9.553756987e-09 wkt1 = -3.972203899e-15 pkt1 = 7.578409011e-22
+ kt2 = -0.028878939
+ at = 5.372048980e+04 lat = -5.378732458e-10 wat = -1.282487996e-09 pat = 2.446807921e-16
+ ute = -1.155115866e+00 lute = -3.064860140e-08 wute = -2.148037751e-07 pute = 4.098155304e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.144 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.145 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.549167264e-01 lvth0 = 5.252285745e-07 wvth0 = -8.881784197e-22
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-07 pk2 = 4.440892099e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.016575863e-01 lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = 3.814697266e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.146 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.031067740e-01 lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-07 pk2 = -1.110223025e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.179965467e-01 lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 2.220446049e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.147 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.427426575e-01 lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.375696972e-01 lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24 pub1 = 3.081487911e-45
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.148 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.911229542e-01 lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.358925766e-02 lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-06 wnfactor = 7.105427358e-21
+ eta0 = -1.553159062e-03 leta0 = 4.128463499e-9
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = 1.561251128e-23 petab = 1.110223025e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = -5.293955920e-29
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = -5.293955920e-28 palpha0 = -5.717472394e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -4.135903063e-31 pua1 = 4.135903063e-37
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 wub1 = -3.851859889e-40 pub1 = -1.540743956e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.149 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.552397824e-01 lvth0 = 1.920515398e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610696e-8
+ k2 = -7.935304322e-02 lk2 = 3.627992986e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667335e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.255026664e-01 lvoff = -9.262472597e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217672e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -2.081668171e-22 peta0 = 2.810252031e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.664850807e-02 lu0 = -4.691369216e-9
+ ua = -6.439244642e-10 lua = -4.848866142e-16
+ ub = 1.111503269e-18 lub = 2.659850321e-25
+ uc = 2.628890915e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111883581e+05 lvsat = 1.967033607e-01 pvsat = -1.164153218e-22
+ a0 = 1.011417809e+00 la0 = 1.906162387e-7
+ ags = 2.367344375e+00 lags = -1.129396051e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608782e-08 lb1 = -3.169227302e-14
+ keta = -1.194413445e-01 lketa = 5.737558585e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701755e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109109e-03 lpdiblc2 = -4.799688220e-9
+ pdiblcb = 9.625889889e-02 lpdiblcb = -9.749071473e-08 wpdiblcb = 4.336808690e-24 ppdiblcb = 2.016616041e-29
+ drout = 8.376749865e-01 ldrout = 8.291329327e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279457e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552343e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457430e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380073e-9
+ at = 1.158432509e+05 lat = -5.372855313e-2
+ ute = -8.338566440e-01 lute = -2.433498184e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563804e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648481e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475369e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.150 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.316084900e-01 lvth0 = -1.980291269e-8
+ k1 = 2.425254334e-02 lk1 = 2.302273434e-7
+ k2 = 1.364915753e-01 lk2 = -7.397047947e-08 wk2 = -8.326672685e-23 pk2 = -2.081668171e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988866e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.072895691e-01 lvoff = -1.856546771e-8
+ nfactor = 4.181852129e+00 lnfactor = -7.003856918e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928472e-02 letab = -2.311014721e-08 wetab = 8.673617380e-24 petab = 2.168404345e-30
+ u0 = 1.451973038e-02 lu0 = 1.503840623e-9
+ ua = -2.102031242e-09 lua = 2.598939142e-16 wua = -3.308722450e-30
+ ub = 2.286030502e-18 lub = -3.339470352e-25
+ uc = 1.078724767e-11 luc = 2.132518899e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.752347497e+05 lvsat = -6.761528150e-4
+ a0 = 1.264221183e+00 la0 = 6.148781451e-8
+ ags = -9.846887499e-01 lags = 5.827755403e-07 wags = -4.440892099e-22 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.220181432e-02 lketa = -4.051305667e-08 wketa = 2.775557562e-23 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500265e-01 lpclm = -1.136192514e-7
+ pdiblc1 = -3.048846468e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = 5.551115123e-29
+ pdiblc2 = -8.673906560e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 3.361026735e-24 ppdiblc2 = -1.978668965e-30
+ pdiblcb = -8.553970447e-02 lpdiblcb = -4.630533306e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076254e+07 lpscbe1 = 1.888714225e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729689e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380753e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373154e+03 lat = 9.625574790e-3
+ ute = -1.301136473e+00 lute = -4.669823687e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393851e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873019e-25 wub1 = 1.540743956e-39
+ uc1 = -1.418079323e-10 luc1 = 7.536563684e-17 wuc1 = -9.047287950e-32 puc1 = 1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.151 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.910376278e-01 lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610978680e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456701426e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016985107e-18
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380979e-02 lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149791621e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.285816312e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026290495e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865197e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.152 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.663494217e-01 lvth0 = 2.487564257e-09 wvth0 = 2.944699932e-08 pvth0 = -5.618075213e-15
+ k1 = 0.90707349
+ k2 = -1.642822690e-02 lk2 = -2.442029014e-08 wk2 = -2.380983222e-08 pk2 = 4.542582650e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.666911915e+00 ldsub = -4.213092735e-07 wdsub = -9.761079297e-07 pdsub = 1.862277275e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079586503e-19
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300002e-01 lvoff = 2.724309667e-17
+ nfactor = -3.997892211e+00 lnfactor = 1.129625373e-06 wnfactor = 1.621326138e-06 pnfactor = -3.093263285e-13
+ eta0 = -1.264693740e-02 leta0 = 2.412858647e-09 weta0 = 3.944984598e-09 peta0 = -7.526478316e-16
+ etab = -0.043998
+ u0 = -1.293558438e-01 lu0 = 2.962168606e-08 wu0 = 5.846163092e-08 pu0 = -1.115366072e-14
+ ua = -1.023245120e-09 lua = -1.325665546e-17 wua = 1.329012897e-16 pua = -2.535570545e-23
+ ub = -4.555562994e-18 lub = 1.140747674e-24 wub = 5.016704073e-25 pub = -9.571169033e-32
+ uc = -2.367505281e-10 luc = 5.985997139e-17 wuc = 1.138127893e-16 puc = -2.171388681e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.842833836e+06 lvsat = -2.962773573e-01 wvsat = -6.372424012e-01 pvsat = 1.215769288e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.404690650e-06 lb0 = -6.525287670e-13 wb0 = -3.644673002e-13 pb0 = 6.953525834e-20
+ b1 = 2.645164180e-06 lb1 = -5.026318756e-13 wb1 = -1.372712398e-12 pb1 = 2.618943076e-19
+ keta = -8.680495464e-01 lketa = 1.604604788e-07 wketa = 3.716866934e-07 pketa = -7.091261748e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.238616222e-02 lpclm = 3.183781848e-08 wpclm = 1.113923637e-07 ppclm = -2.125210350e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000016e-08 lalpha0 = -2.923100113e-23 walpha0 = 2.103028225e-22 palpha0 = -4.012283898e-29
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968489e-08 wbeta0 = 3.808509064e-17 pbeta0 = -7.275957614e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.815416658e-01 lkt1 = -9.553755267e-09 wkt1 = -7.824496606e-17 pkt1 = 1.492805879e-23
+ kt2 = -0.028878939
+ at = 5.372048689e+04 lat = 1.763598993e-11 wat = -2.483697608e-11 pat = 4.738511052e-18
+ ute = -1.159677081e+00 lute = -2.977838545e-08 wute = -2.128336404e-07 pute = 4.060567893e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.153 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.154 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.305913336e-01 lvth0 = 1.011998805e-06 wvth0 = 1.002040773e-08 pvth0 = -2.005162347e-13
+ k1 = 7.868894831e-01 lk1 = -4.379996120e-06 wk1 = -7.182648365e-08 pk1 = 1.437304393e-12
+ k2 = -1.195722482e-01 lk2 = 1.753665286e-06 wk2 = 3.054281727e-08 pk2 = -6.111857802e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.014231969e-01 lvoff = -1.371667962e-07 wvoff = -9.655247898e-11 pvoff = 1.932090995e-15
+ nfactor = 4.776205409e+00 lnfactor = -1.708931949e-05 wnfactor = -1.724151410e-07 pnfactor = 3.450162491e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.586123952e-02 lu0 = 1.229274687e-07 wu0 = 1.508846931e-09 pu0 = -3.019321304e-14
+ ua = -1.567945616e-09 lua = 1.038160210e-14 wua = 1.362153298e-16 pua = -2.725775815e-21
+ ub = 1.305420030e-18 lub = -1.142016165e-24 wub = -5.318277982e-27 pub = 1.064229226e-31
+ uc = 6.333423789e-11 luc = -2.961043608e-16 wuc = 1.458237511e-20 puc = -2.918047878e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.116168035e+00 la0 = 4.931297306e-06 wa0 = 1.132278538e-07 pa0 = -2.265778352e-12
+ ags = 3.189492136e-01 lags = 5.188954170e-07 wags = 7.462744911e-10 pags = -1.493353914e-14
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.577685926e-08 lb0 = -8.020494973e-13 wb0 = -1.548761980e-14 pb0 = 3.099194454e-19
+ b1 = 1.533352558e-08 lb1 = -5.920242223e-14 wb1 = 7.533083426e-16 pb1 = -1.507429204e-20
+ keta = -4.819492937e-03 lketa = 5.460802153e-09 wketa = 8.927844716e-10 pketa = -1.786531901e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.567951267e-02 lpclm = -5.764009390e-07 wpclm = -2.286516418e-08 ppclm = 4.575499072e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 2.763457643e-03 lpdiblc2 = -3.608205223e-08 wpdiblc2 = -9.118428639e-10 ppdiblc2 = 1.824669241e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -1.004485635e+08 lpscbe1 = 6.512481558e+03 wpscbe1 = 1.031667870e+01 ppscbe1 = -2.064448497e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.979454292e-01 lkt1 = 2.314333279e-07 wkt1 = 6.073130341e-09 pkt1 = -1.215281116e-13
+ kt2 = -5.740837429e-02 lkt2 = 5.581096922e-07 wkt2 = 9.028723014e-09 pkt2 = -1.806718441e-13
+ at = 2.296000487e+05 lat = -1.092589891e+00 wat = -1.286680157e-02 pat = 2.574748127e-7
+ ute = -6.770835021e-01 lute = -8.771057639e-06 wute = -1.393903503e-07 pute = 2.789310471e-12
+ ua1 = 1.509250306e-09 lua1 = -7.769193781e-15 wua1 = -1.976340721e-16 pua1 = 3.954813123e-21
+ ub1 = -8.022631173e-19 lub1 = 4.658373252e-24 wub1 = 1.731785713e-25 pub1 = -3.465439329e-30
+ uc1 = 1.513892071e-10 luc1 = -2.352685020e-15 wuc1 = -3.374747090e-17 puc1 = 6.753134183e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.155 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.251093781e-01 lvth0 = 2.548349776e-07 wvth0 = -9.063576713e-09 pvth0 = -4.763851928e-14
+ k1 = -9.731408218e-02 lk1 = 2.703169421e-06 wk1 = 2.198486255e-07 pk1 = -8.992424877e-13
+ k2 = 2.511914443e-01 lk2 = -1.216443311e-06 wk2 = -9.485651157e-08 pk2 = 3.933614077e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.283237652e-02 lvoff = -2.059860198e-07 wvoff = -1.036592696e-08 pvoff = 8.419785228e-14
+ nfactor = 3.799359222e+00 lnfactor = -9.264013724e-06 wnfactor = 8.042150399e-08 pnfactor = 1.424742234e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.111833772e-02 lu0 = 7.061200158e-10 wu0 = -3.050535332e-09 pu0 = 6.331022559e-15
+ ua = -1.238479865e-10 lua = -1.186754974e-15 wua = -3.504206920e-16 pua = 1.172561216e-21
+ ub = 9.800139738e-19 lub = 1.464742117e-24 wub = 1.532480793e-25 pub = -1.163818232e-30
+ uc = -6.280647041e-11 luc = 7.143818593e-16 wuc = 2.976625492e-17 puc = -2.386260867e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.047189575e+00 la0 = -2.526917007e-06 wa0 = -2.623788062e-07 pa0 = 7.431262215e-13
+ ags = 2.172567339e-01 lags = 1.333532110e-06 wags = 5.912826808e-08 pags = -4.826191961e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.729213055e-07 lb0 = 7.896789789e-13 wb0 = 7.069918857e-14 pb0 = -3.805046325e-19
+ b1 = 1.474336057e-08 lb1 = -5.447473666e-14 wb1 = -3.564313932e-15 pb1 = 1.951325603e-20
+ keta = -1.198656708e-02 lketa = 6.287469937e-08 wketa = -2.292473845e-09 pketa = 7.651103722e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.799318387e+00 lpclm = 1.420348241e-05 wpclm = 4.523878342e-07 ppclm = -3.349600158e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -3.516886206e-03 lpdiblc2 = 1.422843835e-08 wpdiblc2 = 7.602127475e-10 ppdiblc2 = 4.852212732e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.915650021e+08 lpscbe1 = -2.235405425e+03 wpscbe1 = -1.453572731e+02 ppscbe1 = 1.040625864e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.975461713e-01 lkt1 = 2.282349584e-07 wkt1 = 4.662816536e-09 pkt1 = -1.102303895e-13
+ kt2 = 1.762431711e-02 lkt2 = -4.296114161e-08 wkt2 = -1.125627331e-08 pkt2 = -1.817307950e-14
+ at = 4.629423130e+04 lat = 3.758337852e-01 wat = 3.860040471e-02 pat = -1.548179628e-7
+ ute = -2.561128647e+00 lute = 6.321624833e-06 wute = 5.480430399e-07 pute = -2.717571307e-12
+ ua1 = -1.235537772e-09 lua1 = 1.421871612e-14 wua1 = 1.134331838e-15 pua1 = -6.715280743e-21
+ ub1 = 1.045270910e-18 lub1 = -1.014182647e-23 wub1 = -8.544585660e-25 pub1 = 4.766741863e-30
+ uc1 = -2.568724225e-10 luc1 = 9.178115262e-16 wuc1 = 7.629790755e-17 puc1 = -2.062365587e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.156 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.449600164e-01 lvth0 = -2.258602848e-07 wvth0 = -4.210660109e-08 pvth0 = 8.488998031e-14
+ k1 = 6.767922676e-01 lk1 = -4.016054889e-07 wk1 = -4.851042420e-08 pk1 = 1.770882319e-13
+ k2 = -1.140809945e-01 lk2 = 2.485862726e-07 wk2 = 2.836213145e-08 pk2 = -1.008422007e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.802460648e+00 ldsub = -4.983243772e-06 wdsub = -3.875632348e-07 pdsub = 1.554433196e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.185389296e-01 lvoff = 2.981960633e-07 wvoff = 3.335381783e-08 pvoff = -9.115268803e-14
+ nfactor = -1.302471700e+00 lnfactor = 1.119833831e-05 wnfactor = 1.308493788e-06 pnfactor = -3.500792888e-12
+ eta0 = 4.092520717e-01 leta0 = -1.320559600e-06 weta0 = -1.027042572e-07 peta0 = 4.119247970e-13
+ etab = -3.578367167e-01 letab = 1.154451474e-06 wetab = 8.978548273e-08 petab = -3.601103571e-13
+ u0 = 3.292302386e-02 lu0 = -6.532089871e-09 wu0 = -1.390777024e-09 pu0 = -3.259128268e-16
+ ua = -1.372457982e-09 lua = 3.821152515e-15 wua = 2.743738166e-16 pua = -1.333355852e-21
+ ub = 3.374251416e-18 lub = -8.138031897e-24 wub = -7.791033910e-25 pub = 2.575643992e-30
+ uc = 1.634440429e-10 luc = -1.930605318e-16 wuc = -5.272783789e-17 puc = 9.224006587e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.932576895e+05 lvsat = -8.553309555e-01 wvsat = -8.784766655e-02 pvsat = 3.523381911e-7
+ a0 = 4.047405694e+00 la0 = -1.054935582e-05 wa0 = -1.001047615e-06 pa0 = 3.705768740e-12
+ ags = -2.910547498e-02 lags = 2.321638208e-06 wags = 1.460667578e-07 pags = -8.313108734e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.094130473e-07 lb0 = 9.360395460e-13 wb0 = 6.545155449e-14 pb0 = -3.594574952e-19
+ b1 = -1.774042840e-08 lb1 = 7.581078938e-14 wb1 = 4.510421413e-15 pb1 = -1.287277944e-20
+ keta = 4.282352676e-02 lketa = -1.569568577e-07 wketa = -1.744319475e-08 pketa = 6.841740302e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.036177216e+00 lpclm = -2.123379966e-05 wpclm = -2.436380297e-06 ppclm = 8.236630620e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.239717606e-02 lpdiblc2 = -4.959945979e-08 wpdiblc2 = -4.104489560e-09 ppdiblc2 = 2.436349264e-14
+ pdiblcb = -7.676919366e-02 lpdiblcb = 2.076351572e-07 wpdiblcb = 1.614846812e-08 ppdiblcb = -6.476804984e-14
+ drout = 0.56
+ pscbe1 = 6.646040177e+07 lpscbe1 = 1.474991155e+03 wpscbe1 = 2.288144740e+02 ppscbe1 = -4.600969408e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.099213957e-01 lkt1 = -5.242878645e-07 wkt1 = -6.102148779e-08 pkt1 = 1.532152987e-13
+ kt2 = 1.182831932e-01 lkt2 = -4.466823525e-07 wkt2 = -5.468480051e-08 pkt2 = 1.560094494e-13
+ at = 2.668552321e+05 lat = -5.087891891e-01 wat = -3.957020627e-02 pat = 1.587076293e-7
+ ute = 1.475554346e+00 lute = -9.868646804e-06 wute = -9.645923141e-07 pute = 3.349285394e-12
+ ua1 = 9.963154521e-09 lua1 = -3.069684215e-14 wua1 = -3.214224497e-15 pua1 = 1.072584813e-20
+ ub1 = -6.397255323e-18 lub1 = 1.970855355e-23 wub1 = 2.017183453e-24 pub1 = -6.750799742e-30
+ uc1 = -1.487316875e-10 luc1 = 4.840821802e-16 wuc1 = 6.456176813e-17 puc1 = -1.591654151e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.157 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.416120062e-01 lvth0 = 1.830290472e-07 wvth0 = 2.039514383e-08 pvth0 = -4.078765335e-14
+ k1 = 4.982244104e-01 lk1 = -4.254374149e-08 wk1 = 3.871683499e-08 pk1 = 1.692880326e-15
+ k2 = 2.288641947e-02 lk2 = -2.682588582e-08 wk2 = -2.723736238e-08 pk2 = 1.095648308e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.621685496e+00 ldsub = 1.901981355e-06 wdsub = 7.751264696e-07 pdsub = -7.834869837e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 4.248839559e-02 lvoff = -2.266740278e-07 wvoff = -4.369677986e-08 pvoff = 6.377957509e-14
+ nfactor = 7.381643048e+00 lnfactor = -6.263558046e-06 wnfactor = -1.300748206e-06 pnfactor = 1.745834383e-12
+ eta0 = -5.001998154e-01 leta0 = 5.081535227e-07 weta0 = 2.054085144e-07 peta0 = -2.076240507e-13
+ etab = 7.852496013e-01 letab = -1.144050491e-06 wetab = -2.887519434e-07 petab = 4.010473998e-13
+ u0 = 3.018844128e-02 lu0 = -1.033429503e-09 wu0 = -1.417053343e-10 pu0 = -2.837528693e-15
+ ua = 1.933638684e-09 lua = -2.826700375e-15 wua = -6.730837394e-16 pua = 5.717785370e-22
+ ub = -2.915551493e-18 lub = 4.509415736e-24 wub = 1.080273374e-24 pub = -1.163164776e-30
+ uc = 1.050319021e-10 luc = -7.560621687e-17 wuc = -1.766516822e-17 puc = 2.173654055e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.805411377e+04 lvsat = -1.489180998e-01 wvsat = 5.544656986e-02 pvsat = 6.420414669e-8
+ a0 = -2.677942814e+00 la0 = 2.973880810e-06 wa0 = 1.303234058e-06 pa0 = -9.276485887e-13
+ ags = -2.303825178e+00 lags = 6.895612740e-06 wags = 8.231973570e-07 pags = -2.192875602e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.447998951e-07 lb0 = 1.811509324e-12 wb0 = 2.423431492e-13 pb0 = -7.151486374e-19
+ b1 = -1.808193556e-08 lb1 = 7.649748719e-14 wb1 = 7.400223458e-15 pb1 = -1.868355294e-20
+ keta = 2.462311287e-01 lketa = -5.659660159e-07 wketa = -7.117456941e-08 pketa = 1.764596990e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.444852107e+00 lpclm = 7.884451368e-06 wpclm = 3.123210116e-06 ppclm = -2.942515948e-12
+ pdiblc1 = 1.167079867e+00 lpdiblc1 = -1.562541318e-06 wpdiblc1 = -3.052679362e-07 ppdiblc1 = 6.138284924e-13
+ pdiblc2 = -2.581068363e-02 lpdiblc2 = 2.722836956e-08 wpdiblc2 = 1.462482297e-08 ppdiblc2 = -1.329714678e-14
+ pdiblcb = -2.475802147e-02 lpdiblcb = 1.030518203e-07 wpdiblcb = -7.548084717e-11 ppdiblcb = -3.214516040e-14
+ drout = -6.406317959e-01 ldrout = 2.414213606e-06 wdrout = 3.448070684e-07 pdrout = -6.933332258e-13
+ pscbe1 = 1.075235807e+09 lpscbe1 = -5.534403071e+02 wpscbe1 = -8.585485570e+01 ppscbe1 = 1.726357419e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.282899291e-05 lalpha0 = 4.596454292e-11 walpha0 = 7.130451377e-12 palpha0 = -1.433781180e-17
+ alpha1 = 0.85
+ beta0 = -1.146158552e+00 lbeta0 = 3.017417353e-05 wbeta0 = 4.680901049e-06 pbeta0 = -9.412290297e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.349159301e-01 lkt1 = 3.302851953e-07 wkt1 = 5.820385706e-08 pkt1 = -8.652135556e-14
+ kt2 = -1.793184377e-01 lkt2 = 1.517308404e-07 wkt2 = 4.518360462e-08 pkt2 = -4.480454149e-14
+ at = 1.766676771e+05 lat = -3.274413161e-01 wat = -8.284856880e-03 pat = 9.579948677e-8
+ ute = -4.694601147e+00 lute = 2.538215479e-06 wute = 9.479945560e-07 pute = -4.965175086e-13
+ ua1 = -9.080467514e-09 lua1 = 7.595806433e-15 wua1 = 3.077194516e-15 pua1 = -1.924849145e-21
+ ub1 = 5.339270394e-18 lub1 = -3.891088049e-24 wub1 = -1.795278181e-24 pub1 = 9.152447362e-31
+ uc1 = 1.641971944e-10 luc1 = -1.451508344e-16 wuc1 = -3.784801648e-17 puc1 = 4.675874607e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.158 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.049961088e-01 lvth0 = 1.788268370e-08 wvth0 = -2.049622307e-08 pvth0 = 5.447678252e-16
+ k1 = 7.571772566e-01 lk1 = -3.042896532e-07 wk1 = -5.028662417e-08 pk1 = 9.165633079e-14
+ k2 = -1.151727407e-01 lk2 = 1.127223804e-07 wk2 = 1.475527961e-08 pk2 = -3.148909155e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.924073019e-01 ldsub = 6.832175295e-08 wdsub = 6.673439569e-09 pdsub = -6.745419288e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -3.146488068e-01 lvoff = 1.343152565e-07 wvoff = 7.791534794e-08 pvoff = -5.914426111e-14
+ nfactor = -4.064411422e+00 lnfactor = 5.305953568e-06 wnfactor = 2.340341541e-06 pnfactor = -1.934528158e-12
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 2.688821388e-23 peta0 = 2.818925648e-29
+ etab = -6.990280776e-01 letab = 3.562366066e-07 wetab = 2.179517475e-07 petab = -1.111215972e-13
+ u0 = 4.827238984e-02 lu0 = -1.931243154e-08 wu0 = -8.907568867e-09 pu0 = 6.022883444e-15
+ ua = 1.278271205e-09 lua = -2.164264102e-15 wua = -7.918139063e-16 pua = 6.917893275e-22
+ ub = -2.326669368e-19 lub = 1.797593587e-24 wub = 5.537067210e-25 pub = -6.309185751e-31
+ uc = -1.459348637e-10 luc = 1.780674764e-16 wuc = 7.094448321e-17 puc = -6.782885457e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.403778985e+05 lvsat = 7.429224293e-01 wvsat = 3.415697057e-01 pvsat = -2.250051133e-7
+ a0 = -5.126263919e-01 la0 = 7.852092845e-07 wa0 = 6.278025757e-07 pa0 = -2.449319025e-13
+ ags = 8.538587052e+00 lags = -4.063745747e-06 wags = -2.542132338e-06 pags = 1.208752539e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.860318738e-06 lb0 = -7.206295186e-13 wb0 = -7.512278901e-13 pb0 = 2.891390592e-19
+ b1 = 1.576279736e-07 lb1 = -1.011076291e-13 wb1 = -3.937323738e-14 pb1 = 2.859440645e-20
+ keta = -6.098014576e-01 lketa = 2.992997378e-07 wketa = 2.019950221e-07 pketa = -9.965629978e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.967141068e-01 lpclm = -4.460083784e-07 wpclm = 2.064539015e-07 ppclm = 5.700398618e-15
+ pdiblc1 = 6.875439659e-01 lpdiblc1 = -1.077833142e-06 wpdiblc1 = -2.021418899e-09 ppdiblc1 = 3.073111581e-13
+ pdiblc2 = 6.305515001e-03 lpdiblc2 = -5.234234385e-09 wpdiblc2 = 1.292475416e-09 ppdiblc2 = 1.790034709e-16
+ pdiblcb = 4.745042074e-01 lpdiblcb = -4.015954510e-07 wpdiblcb = -1.558113464e-07 ppdiblcb = 1.252704722e-13
+ drout = 2.511772333e+00 ldrout = -7.721923531e-07 wdrout = -6.896142680e-07 pdrout = 3.522453791e-13
+ pscbe1 = 1.777321433e+09 lpscbe1 = -1.263098629e+03 wpscbe1 = -3.048578294e+02 ppscbe1 = 3.940008816e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.127868928e-05 lalpha0 = -8.726744729e-12 walpha0 = -9.929102912e-12 palpha0 = 2.905746839e-18
+ alpha1 = 0.85
+ beta0 = 3.191939782e+01 lbeta0 = -3.248027931e-06 wbeta0 = -6.187774215e-06 pbeta0 = 1.573614498e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.214628087e-01 lkt1 = 1.345116850e-08 wkt1 = -2.010601048e-08 pkt1 = -7.366837796e-15
+ kt2 = -6.347895933e-02 lkt2 = 3.464191743e-08 wkt2 = 1.901180946e-08 pkt2 = -1.835045736e-14
+ at = -3.425754759e+05 lat = 1.974023935e-01 wat = 1.888373430e-01 pat = -1.034488731e-7
+ ute = -3.630682652e+00 lute = 1.462821559e-06 wute = 1.152102131e-06 pute = -7.028265880e-13
+ ua1 = -5.458360167e-09 lua1 = 3.934631036e-15 wua1 = 2.965713872e-15 pua1 = -1.812166071e-21
+ ub1 = 5.839485692e-18 lub1 = -4.396698668e-24 wub1 = -2.697808360e-24 pub1 = 1.827509606e-30
+ uc1 = 3.562791845e-10 luc1 = -3.393046209e-16 wuc1 = -1.150227729e-16 puc1 = 1.247659095e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.159 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 7.279779487e-01 lvth0 = -4.493471836e-08 wvth0 = -3.969766388e-08 pvth0 = 1.035259497e-14
+ k1 = -6.163447123e-01 lk1 = 3.972861393e-07 wk1 = 2.638825087e-07 pk1 = -6.881686392e-14
+ k2 = 3.690765777e-01 lk2 = -1.346253919e-07 wk2 = -9.580920520e-08 pk2 = 2.498569939e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.879857035e-01 ldsub = 7.058024352e-08 wdsub = -1.334687914e-08 pdsub = 3.480679223e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 8.056854541e-02 lvoff = -6.755623395e-08 wvoff = -7.738476881e-08 pvoff = 2.018086432e-14
+ nfactor = 1.135890527e+01 lnfactor = -2.572060672e-06 wnfactor = -2.956457855e-06 pnfactor = 7.710028181e-13
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.262765349e-02 letab = -2.259075767e-08 wetab = 8.204166366e-10 petab = -2.139531730e-16
+ u0 = 2.161853998e-04 lu0 = 5.234004905e-09 wu0 = 5.892087891e-09 pu0 = -1.536574033e-15
+ ua = -4.892218647e-09 lua = 9.875357269e-16 wua = 1.149367478e-15 pua = -2.997389472e-22
+ ub = 5.666131430e-18 lub = -1.215430036e-24 wub = -1.392371736e-24 pub = 3.631110555e-31
+ uc = 3.175505559e-10 luc = -5.867438711e-17 wuc = -1.263656231e-16 puc = 3.295438538e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.659573895e+05 lvsat = -1.286497472e-01 wvsat = -2.021443585e-01 pvsat = 5.271641867e-8
+ a0 = 5.287516015e-01 la0 = 2.532879847e-07 wa0 = 3.029634556e-07 pa0 = -7.900862772e-14
+ ags = -1.133500860e-01 lags = 3.555426155e-07 wags = -3.589322785e-07 pags = 9.360451319e-14
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.183809937e-07 lb0 = -2.395009058e-13 wb0 = -3.783105195e-13 pb0 = 9.865808713e-20
+ b1 = -8.237386775e-08 lb1 = 2.148195148e-14 wb1 = 3.393243209e-14 pb1 = -8.849103235e-21
+ keta = 3.802209938e-02 lketa = -3.159946554e-08 wketa = 1.407971833e-08 pketa = -3.671793425e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -4.050947308e-01 lpclm = 1.678587505e-07 wpclm = 4.446166446e-07 ppclm = -1.159497963e-13
+ pdiblc1 = -3.278954597e+00 lpdiblc1 = 9.481987926e-07 wpdiblc1 = 1.225114583e-06 ppdiblc1 = -3.194927315e-13
+ pdiblc2 = -1.682264780e-02 lpdiblc2 = 6.579307378e-09 wpdiblc2 = 3.356727276e-09 ppdiblc2 = -8.753874793e-16
+ pdiblcb = -5.291490169e-01 lpdiblcb = 1.110565648e-07 wpdiblcb = 1.827368713e-07 ppdiblcb = -4.765521772e-14
+ drout = 1.518100973e+00 ldrout = -2.646389342e-07 wdrout = 2.625333235e-13 pdrout = -6.846501532e-20
+ pscbe1 = -2.246635793e+09 lpscbe1 = 7.922823868e+02 wpscbe1 = 9.531350815e+02 ppscbe1 = -2.485642854e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.897735550e-05 lalpha0 = -7.551255653e-12 walpha0 = -8.663599683e-12 palpha0 = 2.259345507e-18
+ alpha1 = 0.85
+ beta0 = 3.728599233e+01 lbeta0 = -5.989209276e-06 wbeta0 = -6.348055768e-06 pbeta0 = 1.655484071e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.473189847e-01 lkt1 = -2.442045880e-08 wkt1 = -7.054682586e-08 pkt1 = 1.839762453e-14
+ kt2 = 3.899590679e-02 lkt2 = -1.770080953e-08 wkt2 = -3.455796499e-08 pkt2 = 9.012233458e-15
+ at = 5.971894237e+04 lat = -8.083963181e-03 wat = -2.797360823e-02 pat = 7.295125396e-9
+ ute = -1.907692392e-01 lute = -2.942380531e-07 wute = -4.573957954e-07 pute = 1.192824199e-13
+ ua1 = 4.611184524e-09 lua1 = -1.208751419e-15 wua1 = -1.189283780e-15 pua1 = 3.101485598e-22
+ ub1 = -6.394172991e-18 lub1 = 1.852082916e-24 wub1 = 1.798027458e-24 pub1 = -4.689003888e-31
+ uc1 = -7.828252591e-10 luc1 = 2.425339814e-16 wuc1 = 2.640555494e-16 puc1 = -6.886199051e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.160 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = -3.179394558e-02 lvth0 = 1.532031549e-07 wvth0 = 2.153710557e-07 pvth0 = -5.616575613e-14
+ k1 = 9.070734895e-01 lk1 = 9.610845453e-17
+ k2 = -2.578321670e-01 lk2 = 2.886363201e-08 wk2 = 4.253156721e-08 pk2 = -1.109163729e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.862269127e+00 ldsub = -3.660494333e-07 wdsub = -5.782038727e-07 pdsub = 1.507874752e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999993e-03 lcdscd = 1.467913464e-18 wcdscd = 7.122653162e-19 pcdscd = -1.857489856e-25
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.930380956e-02 lvoff = -2.064804199e-08 wvoff = -9.330769490e-17 pvoff = 2.433334090e-23
+ nfactor = -1.228664795e+01 lnfactor = 3.594368570e-06 wnfactor = 5.198373782e-06 pnfactor = -1.355663105e-12
+ eta0 = 2.586026044e-03 leta0 = -4.933773123e-10 weta0 = 9.052863693e-16 peta0 = -2.360860111e-22
+ etab = -4.399800002e-02 letab = 4.149736110e-18
+ u0 = -3.673397487e-02 lu0 = 1.487008940e-08 wu0 = 1.717967839e-08 pu0 = -4.480219608e-15
+ ua = -1.206504277e-09 lua = 2.635301933e-17 wua = 2.734282884e-17 pua = -7.130626962e-24
+ ub = -2.283224180e-18 lub = 8.576506162e-25 wub = 8.852617319e-25 pub = -2.308638660e-31
+ uc = 2.578509145e-10 luc = -4.310555642e-17 wuc = -5.062348271e-17 puc = 1.320189556e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.212823632e+04 lvsat = 9.512697086e-02 wvsat = 1.308805311e-01 pvsat = -3.413181018e-8
+ a0 = 1.499999998e+00 la0 = 2.935935939e-16
+ ags = 1.250000000e+00 lags = 6.286082765e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.239601204e-07 lb0 = 1.105628639e-13 wb0 = 1.920701509e-13 pb0 = -5.008920638e-20
+ b1 = -4.775969536e-07 lb1 = 1.245505991e-13 wb1 = 1.848007519e-13 pb1 = -4.819344888e-20
+ keta = -5.879486345e-01 lketa = 1.316449383e-07 wketa = 1.449046846e-07 pketa = -3.778911308e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.162516963e-01 lpclm = -4.633689883e-08 wpclm = -6.607551306e-09 ppclm = 1.723156875e-15
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026246086e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347651157e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662110532e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629947662e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.823435072e-07 lalpha0 = -4.191965620e-14 walpha0 = -7.564629709e-14 palpha0 = 1.972749523e-20
+ alpha1 = 0.85
+ beta0 = 2.012949758e+01 lbeta0 = -1.515035635e-06 wbeta0 = -1.880182208e-06 pbeta0 = 4.903251974e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.758255074e-01 lkt1 = -1.698635676e-08 wkt1 = -3.732126582e-08 pkt1 = 9.732863628e-15
+ kt2 = -2.887893901e-02 lkt2 = 1.595196197e-18
+ at = -1.244348822e+05 lat = 3.994077611e-02 wat = 3.502143379e-02 pat = -9.133099632e-9
+ ute = -1.015837471e+00 lute = -7.907180915e-08 wute = -1.285865742e-07 pute = 3.353357834e-14
+ ua1 = -2.384733758e-11 lua1 = 3.009865455e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190878198e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.161 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 1.239660536e+00 lvth0 = -8.937255989e-08 wvth0 = -2.479113947e-07 pvth0 = 3.222204945e-14
+ k1 = 0.90707349
+ k2 = 6.024711742e-02 lk2 = -3.182144236e-08 wk2 = -5.539486016e-08 pk2 = 7.591354085e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -7.208291699e-01 ldsub = 1.267695583e-07 wdsub = 4.194110310e-07 pdsub = -3.954348187e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000005e-03 lcdscd = -8.566584941e-19 wcdscd = -1.661955296e-18 pcdscd = 2.672189726e-25
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -2.075300007e-01 lvoff = 1.122231197e-16 wvoff = 2.177178438e-16 pvoff = -3.500599810e-23
+ nfactor = 2.544759612e+01 lnfactor = -3.604796918e-06 wnfactor = -1.050821276e-05 pnfactor = 1.640933715e-12
+ eta0 = -1.264693491e-02 leta0 = 2.412858568e-09 weta0 = 3.944984094e-09 peta0 = -7.526477988e-16
+ etab = -0.043998
+ u0 = 1.596124794e-01 lu0 = -2.259006522e-08 wu0 = -6.057366839e-08 pu0 = 1.035403041e-14
+ ua = -8.683663778e-10 lua = -3.815895797e-17 wua = 6.910177977e-17 pua = -1.509765017e-23
+ ub = 4.588753830e-19 lub = 3.344964090e-25 wub = -1.563937222e-24 pub = 2.364090056e-31
+ uc = -5.103733979e-10 luc = 1.034608872e-16 wuc = 2.265268053e-16 puc = -3.967449928e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.098033487e+05 lvsat = -3.879174852e-02 wvsat = -1.293176865e-01 pvsat = 1.551036697e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.492642732e-06 lb0 = -8.274561278e-13 wb0 = -8.126295770e-13 pb0 = 1.415934359e-19
+ b1 = 3.691851968e-06 lb1 = -6.709218828e-13 wb1 = -1.803876592e-12 pb1 = 3.312183469e-19
+ keta = -4.725592225e-02 lketa = 2.848833847e-08 wketa = 3.357553419e-08 pketa = -1.654906979e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.504117521e-02 lpclm = 3.785560295e-08 wpclm = 1.268098817e-07 ppclm = -2.373102149e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.984882588e-07 lalpha0 = 6.889491310e-14 walpha0 = 1.765080257e-13 palpha0 = -2.838001940e-20
+ alpha1 = 0.85
+ beta0 = 3.283486342e+00 lbeta0 = 1.698947464e-06 wbeta0 = 4.387091812e-06 pbeta0 = -7.053829438e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.929429503e-01 lkt1 = 2.443661169e-08 wkt1 = 8.708295386e-08 pkt1 = -1.400171983e-14
+ kt2 = -0.028878939
+ at = 2.520946815e+05 lat = -3.189579323e-02 wat = -8.171667875e-02 pat = 1.313889791e-8
+ ute = -1.912586392e+00 lute = 9.201533043e-08 wute = 9.731379786e-08 pute = -9.565050043e-15
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.162 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.163 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.627150263e-01 lvth0 = 3.691784641e-7
+ k1 = 5.566262089e-01 lk1 = 2.277529835e-7
+ k2 = -2.165726269e-02 lk2 = -2.056905354e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.017327274e-01 lvoff = -1.309728469e-7
+ nfactor = 4.223472310e+00 lnfactor = -6.028695726e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.069834161e-02 lu0 = 2.613325382e-8
+ ua = -1.131262846e-09 lua = 1.643236638e-15
+ ub = 1.288370552e-18 lub = -8.008426962e-25
+ uc = 6.338098646e-11 luc = -2.970398364e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.479156936e+00 la0 = -2.332395909e-6
+ ags = 3.213416405e-01 lags = 4.710210753e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.387376907e-08 lb0 = 1.914986009e-13
+ b1 = 1.774850174e-08 lb1 = -1.075279933e-13
+ keta = -1.957380452e-03 lketa = -5.181231829e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.762224597e-02 lpclm = 8.904248667e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.597527482e-04 lpdiblc2 = 2.241368535e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.737507727e+07 lpscbe1 = 5.850655103e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.784760245e-01 lkt1 = -1.581647627e-7
+ kt2 = -2.846385108e-02 lkt2 = -2.109296763e-8
+ at = 1.883513100e+05 lat = -2.671702072e-01 wat = 1.164153218e-16
+ ute = -1.123944838e+00 lute = 1.709889326e-7
+ ua1 = 8.756696787e-10 lua1 = 4.909252558e-15
+ ub1 = -2.470825931e-19 lub1 = -6.451225409e-24
+ uc1 = 4.320065665e-11 luc1 = -1.877470904e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.164 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.960531199e-01 lvth0 = 1.021141305e-7
+ k1 = 6.074825579e-01 lk1 = -1.796463452e-7
+ k2 = -5.290211314e-02 lk2 = 4.460527524e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.260637441e-01 lvoff = 6.393772087e-8
+ nfactor = 4.057176644e+00 lnfactor = -4.696536728e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.133884946e-02 lu0 = 2.100228251e-8
+ ua = -1.247236071e-09 lua = 2.572273326e-15
+ ub = 1.471300791e-18 lub = -2.266257692e-24
+ uc = 3.261899065e-11 luc = -5.061207102e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.206048537e+00 la0 = -1.445829675e-7
+ ags = 4.068117269e-01 lags = -2.136614964e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.372805585e-08 lb0 = -4.301530117e-13 wb0 = 3.541366997e-30 pb0 = -3.319062208e-35
+ b1 = 3.316787051e-09 lb1 = 8.081384646e-15
+ keta = -1.933584143e-02 lketa = 8.740281358e-08 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.490412944e-01 lpclm = 3.465244080e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -1.079775722e-03 lpdiblc2 = 2.978379250e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.255747443e+08 lpscbe1 = 1.100660974e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.825979885e-01 lkt1 = -1.251445908e-7
+ kt2 = -1.846134680e-02 lkt2 = -1.012208889e-7
+ at = 1.700404475e+05 lat = -1.204858063e-1
+ ute = -8.041975216e-01 lute = -2.390438396e-6
+ ua1 = 2.400933761e-09 lua1 = -7.309311599e-15
+ ub1 = -1.693975356e-18 lub1 = 5.139522876e-24 pub1 = 3.081487911e-45
+ uc1 = -1.227453723e-11 luc1 = 2.566528161e-16 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.165 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.099735415e-01 lvth0 = 4.628229852e-8
+ k1 = 5.212762443e-01 lk1 = 1.661087306e-7
+ k2 = -2.315691021e-02 lk2 = -7.469636824e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.116123628e-01 lvoff = 5.976323031e-9
+ nfactor = 2.892332897e+00 lnfactor = -2.459773863e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.846443345e-02 lu0 = -7.576909981e-9
+ ua = -4.928630170e-10 lua = -4.533555576e-16
+ ub = 8.765807986e-19 lub = 1.190369253e-25
+ uc = -5.592278815e-12 luc = 1.026451536e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.163327600e+04 lvsat = 2.742042995e-1
+ a0 = 8.382203100e-01 la0 = 1.330697336e-6
+ ags = 4.391592679e-01 lags = -3.434005609e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.133074850e-10 lb0 = -2.163189654e-13
+ b1 = -3.280798056e-09 lb1 = 3.454288663e-14
+ keta = -1.309633638e-02 lketa = 6.237749411e-08 wketa = 1.734723476e-24 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.744363068e-01 lpclm = 5.171412440e-06 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -7.611070267e-04 lpdiblc2 = 2.850568056e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.055457235e-01 lkt1 = -3.310613675e-8
+ kt2 = -5.702681193e-02 lkt2 = 5.345693870e-8
+ at = 140000.0
+ ute = -1.616761652e+00 lute = 8.685824428e-7
+ ua1 = -3.410928692e-10 lua1 = 3.688370421e-15
+ ub1 = 6.948567385e-20 lub1 = -1.933341932e-24
+ uc1 = 5.824216620e-11 luc1 = -2.617459078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.166 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.069953072e-01 lvth0 = 5.227089047e-8
+ k1 = 6.223438819e-01 lk1 = -3.711666019e-8
+ k2 = -6.443184982e-02 lk2 = 8.298702475e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.759591720e-02 lvoff = -2.220774955e-8
+ nfactor = 3.211669446e+00 lnfactor = -6.667151992e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -1.404391494e-01 letab = 1.416380554e-7
+ u0 = 2.973415850e-02 lu0 = -1.013005535e-8
+ ua = -2.241512811e-10 lua = -9.936773541e-16
+ ub = 5.476179603e-19 lub = 7.805107952e-25
+ uc = 4.840043040e-11 luc = -5.922630220e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.196979920e+05 lvsat = 5.690928146e-2
+ a0 = 1.5
+ ags = 3.352030625e-01 lags = -1.343668785e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.321102943e-07 lb0 = -4.811334227e-13 pb0 = -1.058791184e-34
+ b1 = 5.641899952e-09 lb1 = 1.660125039e-14
+ keta = 1.805777867e-02 lketa = -2.667642893e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.567618932e+00 lpclm = -1.548745445e-6
+ pdiblc1 = 1.884437022e-01 lpdiblc1 = 4.052865819e-7
+ pdiblc2 = 2.107396742e-02 lpdiblc2 = -1.539998143e-8
+ pdiblcb = -0.025
+ drout = 4.647599830e-01 ldrout = 1.915072929e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.483244388e-01 lkt1 = 5.291270522e-8
+ kt2 = -3.446762206e-02 lkt2 = 8.095235534e-9
+ at = 1.501078600e+05 lat = -2.032474338e-2
+ ute = -1.655494688e+00 lute = 9.464662882e-7
+ ua1 = 7.844854756e-10 lua1 = 1.425073244e-15
+ ub1 = -4.160807111e-19 lub1 = -9.569718432e-25
+ uc1 = 4.286300461e-11 luc1 = 4.749612046e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.167 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.392887653e-01 lvth0 = 1.962911505e-8
+ k1 = 5.959670436e-01 lk1 = -1.045532135e-8
+ k2 = -6.786986822e-02 lk2 = 1.177380334e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.138011941e-01 ldsub = 4.669710627e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.486568763e-02 lvoff = -5.529100738e-8
+ nfactor = 3.438318471e+00 lnfactor = -8.958088615e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 1.214306433e-23 peta0 = 7.372574773e-29
+ etab = -0.0003125
+ u0 = 1.971626586e-02 lu0 = -4.109710889e-12
+ ua = -1.260147125e-09 lua = 5.349274039e-17
+ ub = 1.542420970e-18 lub = -2.250221600e-25
+ uc = 8.150086973e-11 luc = -3.938009089e-17 wuc = -5.169878828e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.546354561e+05 lvsat = 2.159498183e-2
+ a0 = 1.5
+ ags = 3.889507903e-01 lags = -1.886943293e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.479878483e-07 lb0 = 2.063002585e-13
+ b1 = 3.140418965e-08 lb1 = -9.438911366e-15
+ keta = 3.775962016e-02 lketa = -2.018110984e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.458569580e+00 lpclm = -4.277338871e-07 wpclm = -8.881784197e-22
+ pdiblc1 = 6.810636468e-01 lpdiblc1 = -9.264676145e-8
+ pdiblc2 = 1.044896747e-02 lpdiblc2 = -4.660380241e-9
+ pdiblcb = -0.025
+ drout = 3.009883541e-01 ldrout = 3.570453626e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.522960400e-07 lalpha0 = 5.885766851e-13 palpha0 = -1.323488980e-35
+ alpha1 = 0.85
+ beta0 = 1.208246472e+01 lbeta0 = 1.796707776e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.859191982e-01 lkt1 = -1.016563836e-8
+ kt2 = -2.530388930e-03 lkt2 = -2.418647259e-8
+ at = 2.628043600e+05 lat = -1.342367878e-1
+ ute = 6.275736411e-02 lute = -7.903188302e-7
+ ua1 = 4.049205174e-09 lua1 = -1.874859721e-15 pua1 = -8.271806126e-37
+ ub1 = -2.809220949e-18 lub1 = 1.461980805e-24
+ uc1 = -1.246391639e-11 luc1 = 6.067328922e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.168 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 2.303300179e-01 lvth0 = 1.774409178e-07 wvth0 = 1.155346505e-07 pvth0 = -5.901348198e-14
+ k1 = 2.296169368e-01 lk1 = 1.766711843e-07 wk1 = -4.134812492e-16 pk1 = 2.112003905e-22
+ k2 = -3.039964410e-02 lk2 = -7.365462557e-09 wk2 = 2.880021162e-08 pk2 = -1.471074489e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.763704446e+00 ldsub = -7.449717762e-07 wdsub = -5.048639779e-07 pdsub = 2.578774518e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446125e-03 lcdscd = -1.783892587e-09 wcdscd = -3.753421185e-18 pcdscd = 1.917195569e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -4.522962738e-01 lvoff = 1.426031120e-07 wvoff = 8.883281999e-08 pvoff = -4.537456079e-14
+ nfactor = -8.485957432e+00 lnfactor = 5.194944330e-06 wnfactor = 3.233789858e-06 pnfactor = -1.651774586e-12
+ eta0 = 9.936117851e-01 leta0 = -2.572377985e-07 weta0 = 2.122630581e-09 peta0 = -1.084209984e-15
+ etab = 4.525776728e-02 letab = -2.327665454e-08 wetab = -1.785311287e-17 petab = 9.119109981e-24
+ u0 = 2.610173547e-02 lu0 = -3.265718191e-09 wu0 = -2.182443512e-09 pu0 = 1.114761592e-15
+ ua = -1.159362785e-09 lua = 2.013510626e-18 wua = -1.502971652e-17 pua = 7.676968781e-24
+ ub = 2.823582036e-18 lub = -8.794212960e-25 wub = -5.056896180e-25 pub = 2.582991772e-31
+ uc = -9.834907063e-11 luc = 5.248474075e-17 wuc = 3.366779216e-18 puc = -1.719703689e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.922456869e+04 lvsat = 1.410474085e-01 wvsat = 6.149494012e-02 pvsat = -3.141075449e-8
+ a0 = 1.500000004e+00 la0 = -2.288416567e-15 wa0 = -1.263108729e-15 pa0 = 6.451776891e-22
+ ags = -1.264024843e+00 lags = 6.556224824e-07 wags = -2.704426127e-16 pags = 1.381386082e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.842282574e-07 lb0 = 4.291257521e-13 wb0 = 2.151741894e-13 pb0 = -1.099079635e-19
+ b1 = -3.866595414e-07 lb1 = 2.041021896e-13 wb1 = 1.288488708e-13 pb1 = -6.581419934e-20
+ keta = 2.279719492e-01 lketa = -1.173389045e-07 wketa = -4.517171822e-08 pketa = 2.307308126e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.573701524e-01 lpclm = 8.366476370e-08 wpclm = 1.755862486e-07 ppclm = -8.968699758e-14
+ pdiblc1 = 6.485507005e-01 lpdiblc1 = -7.603960369e-08 wpdiblc1 = 2.162416912e-16 ppdiblc1 = -1.104530911e-22
+ pdiblc2 = -6.061561146e-03 lpdiblc2 = 3.772966630e-09 wpdiblc2 = -5.797922906e-18 ppdiblc2 = 2.961499102e-24
+ pdiblcb = 5.667376276e-02 lpdiblcb = -4.171781459e-08 wpdiblcb = -1.716726761e-17 ppdiblcb = 8.768791249e-24
+ drout = 1.518101819e+00 ldrout = -2.646391555e-07 wdrout = -1.145304296e-15 pdrout = 5.850055995e-22
+ pscbe1 = 8.089503011e+08 lpscbe1 = -4.571688497e+00 wpscbe1 = -1.131458282e-07 ppscbe1 = 5.779361725e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.497450161e-06 lalpha0 = -4.584049782e-13 walpha0 = -9.173785118e-14 palpha0 = 4.685841005e-20
+ alpha1 = 0.85
+ beta0 = 1.771947945e+01 lbeta0 = -1.082600432e-06 wbeta0 = -2.446342721e-07 pbeta0 = 1.249557613e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.774161146e-01 lkt1 = -6.558749441e-08 wkt1 = -6.115856793e-08 pkt1 = 3.123894028e-14
+ kt2 = -7.179094734e-02 lkt2 = 1.119085100e-08 wkt2 = -6.862899138e-18 pkt2 = 3.505473689e-24
+ at = 1.170882334e+05 lat = -5.980703039e-02 wat = -4.586892592e-02 pat = 2.342920520e-8
+ ute = -1.264973424e+00 lute = -1.121325321e-07 wute = -1.223171357e-07 pute = 6.247788049e-14
+ ua1 = 7.985465814e-10 lua1 = -2.144688213e-16 wua1 = -1.294916094e-24 pua1 = 6.614250949e-31
+ ub1 = -6.300081721e-19 lub1 = 3.488694277e-25 wub1 = -1.839490838e-33 pub1 = 9.395863253e-40
+ uc1 = 6.369112720e-11 luc1 = 2.177435912e-17 wuc1 = 2.663459534e-26 puc1 = -1.360456199e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.169 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 1.981448708e+00 lvth0 = -2.792263209e-07 wvth0 = -4.126237517e-07 pvth0 = 7.872283510e-14
+ k1 = 9.070734848e-01 lk1 = 9.993081918e-16 wk1 = 1.476717415e-15 pk1 = -2.817370781e-22
+ k2 = 2.082612952e-01 lk2 = -6.960489427e-08 wk2 = -1.028578986e-07 pk2 = 1.962384705e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -5.771732862e+00 ldsub = 1.220164778e-06 wdsub = 1.803085635e-06 pdsub = -3.440034961e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999952e-03 lcdscd = 9.071346105e-18 wcdscd = 1.340508607e-17 pcdscd = -2.557501953e-24
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = 9.177770648e-01 lvoff = -2.146928337e-07 wvoff = -3.172600714e-07 pvoff = 6.052877998e-14
+ nfactor = 4.140333344e+01 lnfactor = -7.815484278e-06 wnfactor = -1.154924949e-05 pnfactor = 2.203435114e-12
+ eta0 = 2.688883937e-02 leta0 = -5.130013596e-09 weta0 = -7.580823504e-09 peta0 = 1.446314993e-15
+ etab = -4.399800023e-02 letab = 4.314765212e-17 wetab = 6.376105199e-17 petab = -1.216469980e-23
+ u0 = -6.646528651e-03 lu0 = 5.274570615e-09 wu0 = 7.794441116e-09 pu0 = -1.487070243e-15
+ ua = -1.290928864e-09 lua = 3.632410216e-17 wua = 5.367755899e-17 pua = -1.024092677e-23
+ ub = -5.235061817e-18 lub = 1.222160200e-24 wub = 1.806034350e-24 pub = -3.445660695e-31
+ uc = 1.341083321e-10 luc = -8.136895467e-18 wuc = -1.202421149e-17 puc = 2.294051213e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.031531142e+06 lvsat = -1.486221303e-01 wvsat = -2.196247862e-01 pvsat = 4.190133445e-8
+ a0 = 1.499999984e+00 la0 = 3.052702979e-15 wa0 = 4.511100826e-15 pa0 = -8.606546587e-22
+ ags = 1.249999997e+00 lags = 6.536122754e-16 wags = 9.658673861e-16 pags = -1.842739294e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.655394992e-06 lb0 = -5.200370366e-13 wb0 = -7.684792480e-13 pb0 = 1.466150818e-19
+ b1 = 1.590082190e-06 lb1 = -3.114043796e-13 wb1 = -4.601745387e-13 pb1 = 8.779485955e-20
+ keta = -6.405975466e-01 lketa = 1.091718600e-07 wketa = 1.613275651e-07 pketa = -3.077904083e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.405423034e+00 lpclm = -4.243601551e-07 wpclm = -6.270937450e-07 ppclm = 1.196407072e-13
+ pdiblc1 = 3.569721527e-01 lpdiblc1 = -5.226161726e-16 wpdiblc1 = -7.722906759e-16 ppdiblc1 = 1.473421385e-22
+ pdiblc2 = 8.406112027e-03 lpdiblc2 = 1.401253419e-17 wpdiblc2 = 2.070686678e-17 ppdiblc2 = -3.950582916e-24
+ pdiblcb = -1.032957702e-01 lpdiblcb = 4.149003363e-17 wpdiblcb = 6.131162245e-17 ppdiblcb = -1.169739305e-23
+ drout = 5.033266455e-01 ldrout = 2.767993390e-15 wdrout = 4.090373373e-15 pdrout = -7.803859781e-22
+ pscbe1 = 7.914198786e+08 lpscbe1 = 2.734546661e-07 wpscbe1 = 4.040946960e-07 ppscbe1 = -7.709574699e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.110507114e-06 lalpha0 = 2.217137678e-13 walpha0 = 3.276351828e-13 palpha0 = -6.250820598e-20
+ alpha1 = 0.85
+ beta0 = 1.130104767e+01 lbeta0 = 5.912367196e-07 wbeta0 = 8.736938288e-07 pbeta0 = -1.666885508e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.956988219e-01 lkt1 = 1.478091797e-07 wkt1 = 2.184234569e-07 pkt1 = -4.167213765e-14
+ kt2 = -2.887893909e-02 lkt2 = 1.658642668e-17 wkt2 = 2.451039371e-17 pkt2 = -4.676245502e-24
+ at = -5.373330741e+05 lat = 1.108568847e-01 wat = 1.638175926e-01 pat = -3.125410322e-8
+ ute = -2.828519362e+00 lute = 2.956183591e-07 wute = 4.368469133e-07 pute = -8.334427521e-14
+ ua1 = -2.384735240e-11 lua1 = 3.129577774e-24 wua1 = 4.624700579e-24 pua1 = -8.823281236e-31
+ ub1 = 7.077531467e-19 lub1 = 4.445715765e-33 wub1 = 6.569610508e-33 pub1 = -1.253389623e-39
+ uc1 = 1.471862503e-10 luc1 = -6.437098847e-26 wuc1 = -9.512349570e-26 puc1 = 1.814823924e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.170 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = -1.307351324e-01 lvth0 = 1.237487853e-07 wvth0 = 1.795588670e-07 pvth0 = -3.425731800e-14
+ k1 = 0.90707349
+ k2 = 9.806228507e-02 lk2 = -4.858046592e-08 wk2 = -6.719062103e-08 pk2 = 1.281902982e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.429490745e+00 ldsub = -5.352998694e-07 wdsub = -8.752065606e-07 pdsub = 1.669771589e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = -1.343760374e+01 lnfactor = 2.647398761e-06 wnfactor = 1.621325400e-06 pnfactor = -3.093261878e-13
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 1.766145641e-01 lu0 = -2.968908023e-08 wu0 = -6.587716269e-08 pu0 = 1.256844036e-14
+ ua = -1.072899214e-09 lua = -5.272902601e-18 wua = 1.329021165e-16 pua = -2.535586320e-23
+ ub = -6.163090404e-18 lub = 1.399215062e-24 wub = 5.016658097e-25 pub = -9.571081316e-32
+ uc = -1.113153575e-10 luc = 3.868650857e-17 wuc = 1.020478326e-16 puc = -1.946929779e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.306845638e+05 lvsat = 7.311235533e-02 wvsat = 1.016641890e-01 pvsat = -1.939610396e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.055917419e-06 lb0 = -5.964511084e-13 wb0 = -3.644689769e-13 pb0 = 6.953557823e-20
+ b1 = 2.309490899e-06 lb1 = -4.486574896e-13 wb1 = -1.372673939e-12 pb1 = 2.618869702e-19
+ keta = -1.131181136e+00 lketa = 2.027683406e-07 wketa = 3.716864939e-07 pketa = -7.091257942e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.438503395e-02 lpclm = 2.990856081e-08 wpclm = 1.113922654e-07 ppclm = -2.125208474e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.673659118e-07 lalpha0 = -2.208651526e-14 walpha0 = 2.542867870e-21 palpha0 = -4.851435998e-28
+ alpha1 = 0.85
+ beta0 = 1.734774328e+01 lbeta0 = -5.623881488e-07 wbeta0 = 1.759190127e-14 pbeta0 = -3.356277034e-21
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.137700705e-01 lkt1 = -2.045047907e-08 wkt1 = -8.760734360e-16 pkt1 = 1.671425220e-22
+ kt2 = -0.028878939
+ at = -9.874845431e+03 lat = 1.022523909e-02 wat = -2.813644242e-10 pat = 5.368038546e-17
+ ute = -9.888383039e-01 lute = -5.536703130e-08 wute = -1.908327907e-07 pute = 3.640822481e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.171 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.481164
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.10827784
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.172 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.627150263e-01 lvth0 = 3.691784641e-7
+ k1 = 5.566262089e-01 lk1 = 2.277529835e-7
+ k2 = -2.165726269e-02 lk2 = -2.056905354e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.017327274e-01 lvoff = -1.309728469e-7
+ nfactor = 4.223472310e+00 lnfactor = -6.028695726e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.069834161e-02 lu0 = 2.613325382e-8
+ ua = -1.131262846e-09 lua = 1.643236638e-15
+ ub = 1.288370552e-18 lub = -8.008426962e-25
+ uc = 6.338098646e-11 luc = -2.970398364e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.479156936e+00 la0 = -2.332395909e-6
+ ags = 3.213416405e-01 lags = 4.710210753e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.387376907e-08 lb0 = 1.914986009e-13
+ b1 = 1.774850174e-08 lb1 = -1.075279933e-13
+ keta = -1.957380452e-03 lketa = -5.181231829e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.762224597e-02 lpclm = 8.904248667e-07 ppclm = -1.110223025e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.597527482e-04 lpdiblc2 = 2.241368535e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.737507727e+07 lpscbe1 = 5.850655103e+03 ppscbe1 = -9.536743164e-19
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.784760245e-01 lkt1 = -1.581647627e-7
+ kt2 = -2.846385108e-02 lkt2 = -2.109296763e-8
+ at = 1.883513100e+05 lat = -2.671702072e-1
+ ute = -1.123944838e+00 lute = 1.709889326e-7
+ ua1 = 8.756696787e-10 lua1 = 4.909252558e-15
+ ub1 = -2.470825931e-19 lub1 = -6.451225409e-24
+ uc1 = 4.320065665e-11 luc1 = -1.877470904e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.173 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 4.960531199e-01 lvth0 = 1.021141305e-7
+ k1 = 6.074825579e-01 lk1 = -1.796463452e-7
+ k2 = -5.290211314e-02 lk2 = 4.460527524e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.260637441e-01 lvoff = 6.393772087e-8
+ nfactor = 4.057176644e+00 lnfactor = -4.696536728e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.133884946e-02 lu0 = 2.100228251e-8
+ ua = -1.247236071e-09 lua = 2.572273326e-15
+ ub = 1.471300791e-18 lub = -2.266257692e-24
+ uc = 3.261899065e-11 luc = -5.061207102e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.206048537e+00 la0 = -1.445829675e-7
+ ags = 4.068117269e-01 lags = -2.136614964e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.372805585e-08 lb0 = -4.301530117e-13 wb0 = -8.530300067e-31 pb0 = 2.874452629e-35
+ b1 = 3.316787051e-09 lb1 = 8.081384646e-15
+ keta = -1.933584143e-02 lketa = 8.740281358e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.490412944e-01 lpclm = 3.465244080e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.079775722e-03 lpdiblc2 = 2.978379250e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.255747443e+08 lpscbe1 = 1.100660974e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.825979885e-01 lkt1 = -1.251445908e-7
+ kt2 = -1.846134680e-02 lkt2 = -1.012208889e-7
+ at = 1.700404475e+05 lat = -1.204858063e-1
+ ute = -8.041975216e-01 lute = -2.390438396e-6
+ ua1 = 2.400933761e-09 lua1 = -7.309311599e-15
+ ub1 = -1.693975356e-18 lub1 = 5.139522876e-24
+ uc1 = -1.227453723e-11 luc1 = 2.566528161e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.174 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.099735415e-01 lvth0 = 4.628229852e-8
+ k1 = 5.212762443e-01 lk1 = 1.661087306e-7
+ k2 = -2.315691021e-02 lk2 = -7.469636824e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.116123628e-01 lvoff = 5.976323031e-9
+ nfactor = 2.892332897e+00 lnfactor = -2.459773863e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.846443345e-02 lu0 = -7.576909981e-9
+ ua = -4.928630170e-10 lua = -4.533555576e-16
+ ub = 8.765807986e-19 lub = 1.190369253e-25
+ uc = -5.592278815e-12 luc = 1.026451536e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.163327600e+04 lvsat = 2.742042995e-1
+ a0 = 8.382203100e-01 la0 = 1.330697336e-6
+ ags = 4.391592679e-01 lags = -3.434005609e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.133074850e-10 lb0 = -2.163189654e-13
+ b1 = -3.280798056e-09 lb1 = 3.454288663e-14
+ keta = -1.309633638e-02 lketa = 6.237749411e-08 wketa = 1.734723476e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.744363068e-01 lpclm = 5.171412440e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -7.611070267e-04 lpdiblc2 = 2.850568056e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.055457235e-01 lkt1 = -3.310613675e-8
+ kt2 = -5.702681193e-02 lkt2 = 5.345693870e-08 wkt2 = -2.775557562e-23
+ at = 140000.0
+ ute = -1.616761652e+00 lute = 8.685824428e-7
+ ua1 = -3.410928692e-10 lua1 = 3.688370421e-15
+ ub1 = 6.948567385e-20 lub1 = -1.933341932e-24
+ uc1 = 5.824216620e-11 luc1 = -2.617459078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.175 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.069953072e-01 lvth0 = 5.227089047e-8
+ k1 = 6.223438819e-01 lk1 = -3.711666019e-8
+ k2 = -6.443184982e-02 lk2 = 8.298702475e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-07 wdsub = -4.440892099e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -9.759591720e-02 lvoff = -2.220774955e-8
+ nfactor = 3.211669446e+00 lnfactor = -6.667151992e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -1.404391494e-01 letab = 1.416380554e-7
+ u0 = 2.973415850e-02 lu0 = -1.013005535e-08 wu0 = -1.387778781e-23
+ ua = -2.241512811e-10 lua = -9.936773541e-16
+ ub = 5.476179603e-19 lub = 7.805107952e-25
+ uc = 4.840043040e-11 luc = -5.922630220e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.196979920e+05 lvsat = 5.690928146e-2
+ a0 = 1.5
+ ags = 3.352030625e-01 lags = -1.343668785e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.321102943e-07 lb0 = -4.811334227e-13 pb0 = -1.058791184e-34
+ b1 = 5.641899952e-09 lb1 = 1.660125039e-14
+ keta = 1.805777867e-02 lketa = -2.667642893e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.567618932e+00 lpclm = -1.548745445e-6
+ pdiblc1 = 1.884437022e-01 lpdiblc1 = 4.052865819e-7
+ pdiblc2 = 2.107396742e-02 lpdiblc2 = -1.539998143e-8
+ pdiblcb = -0.025
+ drout = 4.647599830e-01 ldrout = 1.915072929e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.483244388e-01 lkt1 = 5.291270522e-8
+ kt2 = -3.446762206e-02 lkt2 = 8.095235534e-9
+ at = 1.501078600e+05 lat = -2.032474338e-2
+ ute = -1.655494688e+00 lute = 9.464662882e-7
+ ua1 = 7.844854756e-10 lua1 = 1.425073244e-15
+ ub1 = -4.160807111e-19 lub1 = -9.569718432e-25
+ uc1 = 4.286300461e-11 luc1 = 4.749612046e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.176 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 5.392887653e-01 lvth0 = 1.962911505e-8
+ k1 = 5.959670436e-01 lk1 = -1.045532135e-8
+ k2 = -6.786986822e-02 lk2 = 1.177380334e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.138011941e-01 ldsub = 4.669710627e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -6.486568763e-02 lvoff = -5.529100738e-8
+ nfactor = 3.438318471e+00 lnfactor = -8.958088615e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -1.214306433e-23 peta0 = -7.112366252e-29
+ etab = -0.0003125
+ u0 = 1.971626586e-02 lu0 = -4.109710889e-12
+ ua = -1.260147125e-09 lua = 5.349274039e-17
+ ub = 1.542420970e-18 lub = -2.250221600e-25
+ uc = 8.150086973e-11 luc = -3.938009089e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.546354561e+05 lvsat = 2.159498183e-2
+ a0 = 1.5
+ ags = 3.889507903e-01 lags = -1.886943293e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.479878483e-07 lb0 = 2.063002585e-13
+ b1 = 3.140418965e-08 lb1 = -9.438911366e-15
+ keta = 3.775962016e-02 lketa = -2.018110984e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.458569580e+00 lpclm = -4.277338871e-7
+ pdiblc1 = 6.810636468e-01 lpdiblc1 = -9.264676145e-8
+ pdiblc2 = 1.044896747e-02 lpdiblc2 = -4.660380241e-9
+ pdiblcb = -0.025
+ drout = 3.009883541e-01 ldrout = 3.570453626e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.522960400e-07 lalpha0 = 5.885766851e-13 walpha0 = -5.293955920e-29 palpha0 = 1.058791184e-34
+ alpha1 = 0.85
+ beta0 = 1.208246472e+01 lbeta0 = 1.796707776e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.859191982e-01 lkt1 = -1.016563836e-8
+ kt2 = -2.530388930e-03 lkt2 = -2.418647259e-8
+ at = 2.628043600e+05 lat = -1.342367878e-1
+ ute = 6.275736411e-02 lute = -7.903188302e-7
+ ua1 = 4.049205174e-09 lua1 = -1.874859721e-15
+ ub1 = -2.809220949e-18 lub1 = 1.461980805e-24
+ uc1 = -1.246391639e-11 luc1 = 6.067328922e-17 puc1 = 1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.177 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 6.401261761e-01 lvth0 = -3.187722263e-8
+ k1 = 2.296169353e-01 lk1 = 1.766711851e-7
+ k2 = 7.175339854e-02 lk2 = -5.954380660e-08 pk2 = 6.938893904e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -2.702515522e-02 ldsub = 1.697078339e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446112e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -1.372102957e-01 lvoff = -1.833839441e-8
+ nfactor = 2.984148331e+00 lnfactor = -6.638251119e-7
+ eta0 = 1.001140660e+00 leta0 = -2.610834421e-7
+ etab = 4.525776721e-02 letab = -2.327665451e-08 wetab = 1.517883041e-24 petab = -2.602085214e-30
+ u0 = 1.836070744e-02 lu0 = 6.882905486e-10
+ ua = -1.212672507e-09 lua = 2.924337024e-17
+ ub = 1.029923927e-18 lub = 3.675415476e-26
+ uc = -8.640725765e-11 luc = 4.638502987e-17 wuc = 6.462348536e-33 puc = 8.077935669e-40
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.388951911e+05 lvsat = 2.963488884e-2
+ a0 = 1.5
+ ags = -1.264024844e+00 lags = 6.556224829e-07 wags = -2.081668171e-22 pags = -5.898059818e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.210151797e-07 lb0 = 3.928719698e-14 wb0 = 1.058791184e-28
+ b1 = 7.036155178e-08 lb1 = -2.933778654e-14 wb1 = -1.323488980e-29 pb1 = -6.617444900e-36
+ keta = 6.774991616e-02 lketa = -3.549973317e-08 wketa = -1.387778781e-23 pketa = -2.602085214e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.080166602e+00 lpclm = -2.344509436e-7
+ pdiblc1 = 6.485507013e-01 lpdiblc1 = -7.603960408e-8
+ pdiblc2 = -6.061561167e-03 lpdiblc2 = 3.772966640e-09 ppdiblc2 = 2.168404345e-31
+ pdiblcb = 5.667376270e-02 lpdiblcb = -4.171781455e-8
+ drout = 1.518101815e+00 ldrout = -2.646391535e-7
+ pscbe1 = 8.089503007e+08 lpscbe1 = -4.571688292e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.172060170e-06 lalpha0 = -2.922003258e-13
+ alpha1 = 0.85
+ beta0 = 1.685177280e+01 lbeta0 = -6.393880214e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.943427775e-01 lkt1 = 4.521560804e-8
+ kt2 = -7.179094737e-02 lkt2 = 1.119085101e-8
+ at = -4.560676369e+04 lat = 2.329529640e-2
+ ute = -1.698826749e+00 lute = 1.094736726e-7
+ ua1 = 7.985465768e-10 lua1 = -2.144688189e-16 wua1 = -2.067951531e-31
+ ub1 = -6.300081786e-19 lub1 = 3.488694311e-25 wub1 = 9.629649722e-41 pub1 = -1.203706215e-47
+ uc1 = 6.369112730e-11 luc1 = 2.177435907e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.178 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = 0.517891
+ k1 = 0.90707349
+ k2 = -0.156571
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.62373
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = 0.43867
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 0.021
+ ua = -1.100537e-9
+ ub = 1.17086e-18
+ uc = 9.1459e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 252532.0
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.0366e-8
+ b1 = -4.2136e-8
+ keta = -0.068376
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.18115
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.16e-8
+ alpha1 = 0.85
+ beta0 = 14.4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 43720.487
+ ute = -1.2790432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.179 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8__vth0_slope_spectre)
+ vth0 = -5.540233200e-01 lvth0 = 2.045062455e-07 wvth0 = 2.988973523e-07 pvth0 = -5.702543026e-14
+ k1 = 0.90707349
+ k2 = -2.325260563e-01 lk2 = 1.449116137e-08 wk2 = 2.601281122e-08 pk2 = -4.962880202e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.308003241e+00 ldsub = -5.121217546e-07 wdsub = -8.409553457e-07 pdsub = 1.604425066e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
*(mismatch parameter sky130_fd_pr__nfet_01v8__voff_slope_spectre)
+ voff = -0.20753
+ nfactor = -1.343760560e+01 lnfactor = 2.647399117e-06 wnfactor = 1.621325926e-06 pnfactor = -3.093262881e-13
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = -1.159522987e-02 lu0 = 6.218713526e-09 wu0 = -1.281479905e-08 pu0 = 2.444884252e-15
+ ua = -1.072897415e-09 lua = -5.273245830e-18 wua = 1.329016093e-16 pua = -2.535576643e-23
+ ub = -6.163134324e-18 lub = 1.399223441e-24 wub = 5.016781923e-25 pub = -9.571317560e-32
+ uc = -9.715009267e-11 luc = 3.598397435e-17 wuc = 9.805419118e-17 puc = -1.870736692e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.616972904e+05 lvsat = -7.806300910e-02 wvsat = -1.217336119e-01 pvsat = 2.322506889e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.055925333e-06 lb0 = -5.964526183e-13 wb0 = -3.644712082e-13 pb0 = 6.953600393e-20
+ b1 = 2.309501807e-06 lb1 = -4.486595707e-13 wb1 = -1.372677015e-12 pb1 = 2.618875569e-19
+ keta = -1.131181040e+00 lketa = 2.027683223e-07 wketa = 3.716864668e-07 pketa = -7.091257426e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.438497216e-02 lpclm = 2.990857260e-08 wpclm = 1.113922828e-07 ppclm = -2.125208807e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.673659202e-07 lalpha0 = -2.208651686e-14 walpha0 = 1.811849002e-22 palpha0 = -3.456754693e-29
+ alpha1 = 0.85
+ beta0 = 1.734774334e+01 lbeta0 = -5.623881607e-07 wbeta0 = 3.171862772e-17 pbeta0 = -6.053824109e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.137700734e-01 lkt1 = -2.045047852e-08 wkt1 = -6.743006153e-17 pkt1 = 1.286470930e-23
+ kt2 = -0.028878939
+ at = -9.874846353e+03 lat = 1.022523927e-02 wat = -2.139387652e-11 pat = 4.081666702e-18
+ ute = -1.015327828e+00 lute = -5.031320101e-08 wute = -1.833645463e-07 pute = 3.498338833e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.047954
+ k1 = 0.43448553
+ k2 = 0.022159346
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.6628421e-10
+ ub = 1.06194446e-18
+ uc = -6.6549964e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011074
+ a0 = 1.198023
+ keta = 0.0051290095
+ a1 = 0.0
+ a2 = 0.9995
+ ags = 0.2608008
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29454245
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.5294758
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0015228006
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1181082000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4485
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.047954
+ k1 = 0.43448553
+ k2 = 0.022159346
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.6628421e-10
+ ub = 1.06194446e-18
+ uc = -6.6549964e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011074
+ a0 = 1.198023
+ keta = 0.0051290095
+ a1 = 0.0
+ a2 = 0.9995
+ ags = 0.2608008
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29454245
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.5294758
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0015228006
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1181082000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4485
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.052801912332 lvth0 = 3.8751001864043e-8
+ k1 = 0.438102126509735 lk1 = -2.89086783119324e-8
+ k2 = 0.021293418608066 lk2 = 6.92165032718695e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 267009.4996875 lvsat = -0.852865182088082
+ ua = -5.79776770650915e-10 lua = 1.07850597768264e-16
+ ub = 1.0476535911495e-18 lub = 1.14231745035677e-25
+ uc = -7.3167975313894e-11 luc = 5.29000013197789e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0108535677424 lu0 = 1.76198954109988e-9
+ a0 = 1.249119756379 la0 = -4.08433644441004e-7
+ keta = 0.0213163689759253 lketa = -1.29391035618573e-07 pketa = 5.04870979341448e-29
+ a1 = 0.0
+ a2 = 1.19866773275 la2 = -1.59201500656442e-6
+ ags = 0.22509732334312 lags = 2.85389956693552e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.306872589892495 lvoff = 9.85589757479963e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.44269527408715 lnfactor = 6.9366607543917e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.429857606134414 lpclm = 3.44816939760565e-06 wpclm = 1.75362289861242e-22 ppclm = -1.40101696767252e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00576487163879899 lpdiblc2 = -2.2394337483051e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01351357083584e-08 lpscbe2 = -6.06727053633572e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.2565334854499 lbeta0 = 1.11096776216837e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.4402431089145e-11 lagidl = 1.24676640282756e-16
+ bgidl = 1361862407.929 lbgidl = -1445.03890435438
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43171925495647 lkt1 = -1.3413416702476e-7
+ kt2 = 0.0096543549776395 lkt2 = -1.37684887171055e-7
+ at = 87886.257761435 lat = 0.0240898603577266
+ ute = -0.47326335220418 lute = 1.06889595266106e-6
+ ua1 = 1.22719499268165e-09 lua1 = 3.06308714678805e-15
+ ub1 = -3.0164578823216e-19 lub1 = -2.07230654258392e-24
+ uc1 = -8.847741670786e-11 luc1 = -1.60686742927228e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.053297910546 lvth0 = 4.07316903799433e-8
+ k1 = 0.42438480066725 lk1 = 2.58692402332454e-8
+ k2 = 0.025136931386954 lk2 = -8.42679530623213e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53437.5
+ ua = -2.3668488550515e-10 lua = -1.26223126467596e-15
+ ub = 9.3695022895943e-19 lub = 5.56307687997067e-25
+ uc = -8.0533404316558e-11 luc = 8.2312648842419e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0129883399648 lu0 = -6.76287749595451e-9
+ a0 = 1.168811571436 la0 = -8.77359177970925e-8
+ keta = -0.005560794812944 lketa = -2.20614361282578e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.09661181618599 lags = 7.98476014873391e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.28931502304321 lvoff = 2.84456768612062e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.6600217141216 lnfactor = -1.74191855955121e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.139268495071432 letab = 2.76612513571563e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.46408247994329 lpclm = -1.21635517851718e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.853824413469e-05 lpdiblc2 = 7.00772972043594e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800438663.92697 lpscbe1 = -1.75173332879876
+ pscbe2 = 8.2920612364473e-09 lpscbe2 = 1.29274878917682e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.9316215559846 lbeta0 = 8.41382277627077e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.3119513782171e-10 lagidl = -6.21824536352518e-17
+ bgidl = 918666228.2536 lbgidl = 324.793241398225
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.46634935213621 lkt1 = 4.15551598678871e-9
+ kt2 = -0.005808862085711 lkt2 = -7.5935034869729e-8
+ at = 106814.086142966 lat = -0.0514953559757196
+ ute = -0.17622069800093 lute = -1.17295765989642e-7
+ ua1 = 2.3392527360435e-09 lua1 = -1.37773529797308e-15
+ ub1 = -1.02790864263458e-18 lub1 = 8.27906511889728e-25
+ uc1 = -2.40574104777601e-10 luc1 = 4.46686741215816e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.046167775834 lvth0 = 2.65189219133937e-8
+ k1 = 0.3573341256955 lk1 = 1.59523898580084e-7
+ k2 = 0.052817427422536 lk2 = -6.36033799128071e-08 wk2 = -5.29395592033938e-23 pk2 = -5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35743.666875 lvsat = 0.0352697899337212
+ ua = -7.6259585024292e-10 lua = -2.13912954047498e-16
+ ub = 1.15066129181608e-18 lub = 1.30309305384519e-25
+ uc = -4.286074864569e-11 luc = 7.21831273276241e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0100904809916 lu0 = -9.86465086033959e-10
+ a0 = 1.282774495506 la0 = -3.1490254493694e-7
+ keta = -0.007016124315302 lketa = -1.91604725286866e-8
+ a1 = 0.0
+ a2 = 0.7006662 la2 = 1.980058382244e-7
+ ags = 0.3794348864849 lags = 2.34714041569902e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.2758638558486 lvoff = 1.6329541478367e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.3656263388154 lnfactor = 4.12637632666988e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.485738951 leta0 = 9.69238578108438e-07 weta0 = -1.32348898008484e-23 peta0 = 2.17725609840999e-28
+ etab = 7.38760593753566 letab = -1.47269923141726e-05 wetab = 1.79663629046518e-21 petab = -5.41158580981614e-28
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.19003522874366 lpclm = 4.2463328176005e-7
+ pdiblc1 = 0.40797495771238 lpdiblc1 = -3.58301662564802e-8
+ pdiblc2 = 0.00023668464555664 lpdiblc2 = 1.92027487552058e-10
+ pdiblcb = -0.0490937606993659 lpdiblcb = 4.80270087649527e-8
+ drout = 0.40544946099372 ldrout = 3.080714623217e-7
+ pscbe1 = 799122672.14606 lpscbe1 = 0.871483095777194
+ pscbe2 = 8.9456362956796e-09 lpscbe2 = -1.00472122431867e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.4349697107106e-05 lalpha0 = 8.84041358658845e-11 walpha0 = -4.73671530539957e-27 palpha0 = -1.36295278593662e-32
+ alpha1 = 1.993338e-10 lalpha1 = -1.980058382244e-16
+ beta0 = -13.444963104552 lbeta0 = 4.30512292903355e-05 pbeta0 = 2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 807380539.7004 lbgidl = 546.623233247484
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.45647670127916 lkt1 = -1.55240141273016e-8
+ kt2 = -0.040468941952306 lkt2 = -6.84578058861025e-9
+ at = 71198.873273608 lat = 0.0194978012148608
+ ute = -0.16704404204188 lute = -1.35587943025743e-7
+ ua1 = 1.4237427767252e-09 lua1 = 4.47185493314543e-16
+ ub1 = -2.9305679836e-20 lub1 = -1.16264672076927e-24
+ uc1 = -2.1433991940186e-11 luc1 = 9.86642697270848e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.5 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.03759870481 lvth0 = 1.8006938040556e-8
+ k1 = 0.55990344532888 lk1 = -4.16959042458991e-8
+ k2 = -0.032308223178728 lk2 = 2.09551636041513e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 45098.15262 lvsat = 0.0259776237727545
+ ua = -6.248841862818e-10 lua = -3.50707182903309e-16
+ ub = 1.10184261276184e-18 lub = 1.788027543989e-25
+ uc = -5.7784011063288e-11 luc = 2.20421563761344e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0109374520724 lu0 = -1.82779364549367e-9
+ a0 = 1.02077705376 la0 = -5.46505301478509e-8
+ keta = -0.0421967749919 lketa = 1.5785804653104e-8
+ a1 = 0.0
+ a2 = 0.9986676 la2 = -9.80102764488e-8
+ ags = 0.39549313889684 lags = 2.18762769235531e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.25992961562244 lvoff = -1.41951321699368e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.9044637782592 lnfactor = -1.22610071755237e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -14.7771435475356 letab = 7.29009560982912e-6
+ dsub = 0.22117665755564 ldsub = 3.85647013369957e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.61200232157372 lpclm = 5.47733370242402e-9
+ pdiblc1 = 0.700518612109228 lpdiblc1 = -3.26424894827736e-7
+ pdiblc2 = 0.00043
+ pdiblcb = 0.220522721398732 lpdiblcb = -2.19793288329408e-07 wpdiblcb = -7.61006163548785e-23 ppdiblcb = 3.47098798297245e-29
+ drout = 0.43496363801256 ldrout = 2.7875390875016e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.7277890069796e-09 lpscbe2 = 2.06348777819499e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.8699694214212e-05 lalpha0 = -4.37588804104509e-11
+ alpha1 = -9.86676e-11 lalpha1 = 9.80102764488e-17
+ beta0 = 50.1127373244192 lbeta0 = -2.00830497383779e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1694552658.6996 lbgidl = -334.638545094944
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43623405628508 lkt1 = -3.56318026204314e-8
+ kt2 = -0.03963756181126 lkt2 = -7.67162207515662e-9
+ at = 106443.99518944 lat = -0.015512517698768
+ ute = -0.23772148631908 lute = -6.53813518823178e-8
+ ua1 = 3.2739786116024e-09 lua1 = -1.39072407043071e-15
+ ub1 = -2.7909917868124e-18 lub1 = 1.58064103336246e-24 pub1 = 1.40129846432482e-45
+ uc1 = -4.6845503746344e-11 luc1 = 3.51086472872139e-17 puc1 = -1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.6 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.990407688308 lvth0 = -5.274183658508e-9
+ k1 = 0.13549433046384 lk1 = 1.6768123966339e-7
+ k2 = 0.11917144163576 lk2 = -5.37755112760986e-08 wk2 = -5.29395592033938e-23 pk2 = -6.31088724176809e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 98492.4114752 lvsat = -0.000363793102352225
+ ua = -6.323516860368e-10 lua = -3.47023181509177e-16
+ ub = 1.1234768802288e-18 lub = 1.68129748155284e-25
+ uc = -2.5953323664251e-11 luc = 6.33886871606827e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01030450598072 lu0 = -1.51553728651644e-9
+ a0 = 1.15780283375864 la0 = -1.2225055440082e-7
+ keta = 0.059635137695792 lketa = -3.44517474884166e-08 wketa = -2.64697796016969e-23
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.33838723259592 lags = 5.80813843947026e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.22035128023192 lvoff = -3.37206289948251e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.1039853562544 lnfactor = 2.72296351999767e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.965309351859001 leta0 = -2.34488165027416e-7
+ etab = 0.0047760499229952 letab = -2.38704054191061e-09 wetab = 2.68833699079734e-24 petab = -1.08468374467889e-30
+ dsub = 0.1852103104408 ldsub = 5.63082670899366e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.47758274175056 lpclm = 7.17916203732222e-8
+ pdiblc1 = -0.334384403489576 lpdiblc1 = 1.84132089081746e-07 wpdiblc1 = 2.11758236813575e-22 ppdiblc1 = 7.57306469012171e-29
+ pdiblc2 = -0.008973522524736 lpdiblc2 = 4.63911499530821e-09 wpdiblc2 = -4.96308367531817e-24 ppdiblc2 = -1.57772181044202e-30
+ pdiblcb = -0.3710028 lpdiblcb = 7.20287293464e-08 wpdiblcb = -4.2351647362715e-22
+ drout = 1.51703456660792 ldrout = -2.55072799021218e-7
+ pscbe1 = 800003445.66608 lpscbe1 = -0.00169987801257321
+ pscbe2 = 9.40358177202e-09 lpscbe2 = -1.27045473300003e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.72393234514e-09 lalpha0 = 3.85984313528668e-15 walpha0 = -3.15544362088405e-30 palpha0 = -2.49204802374325e-36
+ alpha1 = 1.973352e-10 lalpha1 = -4.80191528976e-17
+ beta0 = 3.3812716986096 lbeta0 = 2.97135805052774e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 484651822.7312 lbgidl = 262.251513520035
+ cgidl = 527.777841138384 lcgidl = -0.000112371464591528
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.45936412512 lkt1 = -2.42208607215494e-8
+ kt2 = 0.00980465974399998 lkt2 = -3.20633487727855e-08 pkt2 = -2.52435489670724e-29
+ at = 63319.776 lat = 0.005762298347712
+ ute = -0.377306802 lute = 3.481388585076e-9
+ ua1 = 7.667833132e-10 lua1 = -1.53829356307462e-16 wua1 = 7.88860905221012e-31 pua1 = 1.88079096131566e-37
+ ub1 = 4.3271957856e-19 lub1 = -9.73828420763331e-27
+ uc1 = 1.101914492e-11 luc1 = 6.56181724345704e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.790897759485714 lvth0 = -5.38225307182653e-8
+ k1 = 0.335246697368572 lk1 = 1.19073898205527e-7
+ k2 = 0.0606923753943428 lk2 = -3.95453322550446e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 158397.929237143 lvsat = -0.0149410819835079
+ ua = -1.56074952462286e-09 lua = -1.21108708263323e-16
+ ub = 1.39430136593714e-18 lub = 1.02227859451988e-25
+ uc = -4.91771559457713e-14 luc = 3.54055130302881e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00571223023114286 lu0 = -3.9806209016584e-10
+ a0 = 0.962178920290572 la0 = -7.46478225453271e-8
+ keta = -0.226972829022943 lketa = 3.52908619169869e-8
+ a1 = 0.0
+ a2 = 0.870068692128286 la2 = -1.70503754051129e-8
+ ags = 4.02569816488 lags = -4.81133968503969e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.149163822694 lvoff = -5.10432425371874e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.604458806285715 lnfactor = 3.93850143616047e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.417167463843577 leta0 = 1.01920978352018e-07 weta0 = -1.12496563307212e-22
+ etab = 0.124203059314531 letab = -3.14481701532282e-08 petab = 3.15544362088405e-30
+ dsub = 0.747409855918 ldsub = -8.04962459073943e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.10997007392457 lpclm = -8.20922482633373e-8
+ pdiblc1 = 1.00596961163057 lpdiblc1 = -1.4202697624956e-07 wpdiblc1 = 1.6940658945086e-21
+ pdiblc2 = 0.0247436758567886 lpdiblc2 = -3.56556062445522e-9
+ pdiblcb = -0.075
+ drout = -0.722076222894571 ldrout = 2.89787942274739e-7
+ pscbe1 = 799987694.049715 lpscbe1 = 0.00213308881063767
+ pscbe2 = 8.09092591147142e-09 lpscbe2 = 1.92373578494165e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.80426155183571e-08 lalpha0 = -4.84351708872099e-15
+ alpha1 = -2.47625714285714e-10 lalpha1 = 6.02567460628571e-17
+ beta0 = 32.89328272192 lbeta0 = -4.21003568786257e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.77947653402857e-11 lagidl = 7.83675739162556e-18
+ bgidl = 2954967410.85428 lbgidl = -338.87014106266
+ cgidl = -513.492289779943 lcgidl = 0.000141009126525876 wcgidl = -2.16840434497101e-19
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.5589
+ kt2 = -0.12196
+ at = 208336.6 lat = -0.0295258055708
+ ute = -0.5190042 lute = 3.79617500196e-8
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.8 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.711113737733333 lvth0 = -6.76521334807794e-8
+ k1 = -0.249508425106668 lk1 = 2.20434181625139e-7
+ k2 = 0.343856885470667 lk2 = -8.86285021026544e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 197157.557086667 lvsat = -0.0216595983556886
+ ua = -9.60007983346665e-10 lua = -2.25240045545056e-16
+ ub = 6.24599095426667e-19 lub = 2.35646511617732e-25
+ uc = 2.69835080537333e-13 luc = -1.98914300172203e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00603241996793333 lu0 = -4.53563138761628e-10
+ a0 = -0.791160669612 la0 = 2.29272555289205e-7
+ keta = -0.0915648642361733 lketa = 1.18195161167778e-8
+ a1 = 0.0
+ a2 = -0.316691314966 la2 = 1.88660230704597e-7
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.390263853465334 lvoff = -9.25144540334603e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -0.669046547333334 lnfactor = 6.14597014601666e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.617243906024667 leta0 = 1.36601828686804e-7
+ etab = -0.246957641957333 letab = 3.28880834838343e-8
+ dsub = 0.393013456590667 ldsub = -1.9065882840793e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.11806085162867 lpclm = -2.5683268748901e-07 wpclm = 3.3881317890172e-21
+ pdiblc1 = 0.985023109708667 lpdiblc1 = -1.38396151499421e-7
+ pdiblc2 = 0.0220607773736267 lpdiblc2 = -3.1005123671809e-9
+ pdiblcb = -0.418610236790253 lpdiblcb = 5.95607112247489e-8
+ drout = 0.709556465021333 ldrout = 4.16315954167721e-8
+ pscbe1 = 867303832.327334 lpscbe1 = -11.6663116879553
+ pscbe2 = 1.013312288888e-08 lpscbe2 = -1.61616761175883e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 14.4732975792 lbeta0 = -1.01715230319377e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.75145547539333e-10 lagidl = -1.0771212493193e-17
+ bgidl = 780957079.713333 lbgidl = 37.9684617166503
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.0674870599999995 lkt1 = -1.0857668020628e-7
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.9 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.062648749802 wvth0 = 1.03594197797603e-7
+ k1 = 0.444388049205489 wk1 = -6.98102075292465e-8
+ k2 = 0.0180906853887137 wk2 = 2.86830084088628e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.9463144281392e-10 wua = 1.99840683421517e-16
+ ub = 1.01974565808793e-18 wub = 2.97490674628997e-25
+ uc = -7.49378332315679e-11 wuc = 5.91323156898652e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01117524733111 wu0 = -7.13767582763556e-10
+ a0 = 1.2066858327441 wa0 = -6.10707375676198e-8
+ keta = 0.0303539152578079 wketa = -1.77829082611841e-7
+ a1 = 0.0
+ a2 = 1.22604688730313 wa2 = -1.59709715169954e-6
+ ags = 0.343036381949931 wags = -5.79739652413986e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.306629209945388 wvoff = 8.52085416482716e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.06134045929744 wnfactor = 3.30023346666222e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.56849442030249 wpclm = 4.018474456923e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0100191156662281 wpdiblc2 = -4.9742059323811e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01311090249299e-08 wpscbe2 = -5.32265564308848e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.342093011489364 wbeta0 = 3.03442588485037e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 268797089.07066 wbgidl = 6431.37343500181
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.479925454664196 wkt1 = 2.21541353900369e-7
+ kt2 = 0.100910653452993 wkt2 = -7.64764870376458e-7
+ at = 93172.3839899999 wat = -0.0160197213089073
+ ute = -0.780957886934979 wute = 3.11188230536035e-6
+ ua1 = 7.2932880804441e-10 wua1 = 6.21132476313363e-15
+ ub1 = -7.73186088509244e-20 wub1 = -3.40912414031835e-24
+ uc1 = -6.65340992675926e-10 wuc1 = 3.92502146538137e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.10 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.062648749802 wvth0 = 1.03594197797603e-7
+ k1 = 0.444388049205489 wk1 = -6.98102075292448e-8
+ k2 = 0.0180906853887137 wk2 = 2.86830084088628e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.94631442813919e-10 wua = 1.99840683421519e-16
+ ub = 1.01974565808792e-18 wub = 2.97490674628997e-25
+ uc = -7.49378332315677e-11 wuc = 5.91323156898654e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01117524733111 wu0 = -7.13767582763556e-10
+ a0 = 1.2066858327441 wa0 = -6.10707375676232e-8
+ keta = 0.0303539152578079 wketa = -1.77829082611841e-7
+ a1 = 0.0
+ a2 = 1.22604688730313 wa2 = -1.59709715169953e-6
+ ags = 0.343036381949931 wags = -5.79739652413987e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.306629209945388 wvoff = 8.52085416482716e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.06134045929744 wnfactor = 3.30023346666222e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.56849442030249 wpclm = 4.018474456923e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0100191156662281 wpdiblc2 = -4.9742059323811e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01311090249299e-08 wpscbe2 = -5.32265564308848e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.342093011489364 wbeta0 = 3.03442588485036e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 268797089.070658 wbgidl = 6431.37343500181
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.479925454664195 wkt1 = 2.21541353900371e-7
+ kt2 = 0.100910653452993 wkt2 = -7.64764870376458e-7
+ at = 93172.3839899999 wat = -0.0160197213089077
+ ute = -0.780957886934979 wute = 3.11188230536035e-6
+ ua1 = 7.29328808044408e-10 wua1 = 6.21132476313363e-15
+ ub1 = -7.73186088509237e-20 wub1 = -3.40912414031835e-24
+ uc1 = -6.65340992675926e-10 wuc1 = 3.92502146538137e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.11 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.06298214945842 lvth0 = 2.66497614281229e-09 wvth0 = 7.17680472761011e-08 pvth0 = 2.5439717835725e-13
+ k1 = 0.417739211580813 lk1 = 2.13013166441158e-07 wk1 = 1.43553300689437e-07 pk1 = -1.70548663805771e-12
+ k2 = 0.0275206297122963 lk2 = -7.53767322995775e-08 wk2 = -4.39002329098013e-08 pk2 = 5.80182380995648e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 275393.831959135 lvsat = -0.919883983839571 wvsat = -0.0591073810341687 pvsat = 4.72465274900901e-7
+ ua = -2.51490382696535e-10 lua = -2.74284247519658e-15 wua = -2.31433440284757e-15 pua = 2.0096651255728e-20
+ ub = 7.43366684165797e-19 lub = 2.20919055465276e-24 wub = 2.14514424907052e-24 pub = -1.47689195274193e-29
+ uc = -9.31427811835541e-11 luc = 1.45518302252635e-16 wuc = 1.40817231876151e-16 puc = -6.52935144578655e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01215566032122 lu0 = -7.83677240953952e-09 wu0 = -9.17941700121389e-09 pu0 = 6.76687971911769e-14
+ a0 = 1.35606158915781 la0 = -1.19401091002048e-06 wa0 = -7.53912351486146e-07 pa0 = 5.53811720051629e-12
+ keta = 0.0733454834213588 lketa = -3.43646135481302e-07 wketa = -3.66791843734603e-07 pketa = 1.51044321906749e-12
+ a1 = 0.0
+ a2 = 1.65138419351546 la2 = -3.39986485256465e-06 wa2 = -3.19153433809292e-06 pa2 = 1.27448753506113e-11
+ ags = 0.418601350570406 lags = -6.0401633514285e-07 wags = -1.36415350661415e-06 pags = 6.27008506850459e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.347588216412412 lvoff = 3.27399182835104e-07 wvoff = 2.87034670476895e-07 pvoff = -1.61326446495874e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.583466011452519 lnfactor = 3.81981198318783e-06 wnfactor = 6.05734479227026e-06 pnfactor = -2.20385227292131e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.55231284286998 lpclm = 7.86399318220881e-06 wpclm = 7.91302005002574e-06 ppclm = -3.11304192820806e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.019740218572311 lpdiblc2 = -7.77040612611031e-08 wpdiblc2 = -9.85225930368203e-08 ppdiblc2 = 3.89919293788478e-13
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.37853598461252e-08 lpscbe2 = -2.92096619505918e-14 wpscbe2 = -2.57331391434733e-14 ppscbe2 = 1.63147893361998e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -3.75323786342985 lbeta0 = 3.27353639050649e-05 wbeta0 = 4.94170808905484e-05 pbeta0 = -1.52455513195914e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.50205801158688e-11 lagidl = 4.39469086177782e-16 wagidl = 2.77631896720417e-16 pagidl = -2.21920559006739e-21
+ bgidl = 765453235.265036 lbgidl = -3969.94044630906 wbgidl = 4204.53091299624 pbgidl = 0.017799904951163
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.488364753628569 lkt1 = 6.74581691052819e-08 wkt1 = 3.99336162428739e-07 pkt1 = -1.42117399921254e-12
+ kt2 = 0.159378129288713 lkt2 = -4.67350296361748e-07 wkt2 = -1.05551401010405e-06 pkt2 = 2.3240561470519e-12
+ at = 93442.9686279172 lat = -0.00216287446848007 wat = -0.0391733790886386 pat = 1.85075012569723e-7
+ ute = -1.35535786977856 lute = 4.59137321006297e-06 wute = 6.21853894493278e-06 pute = -2.48325565700466e-11
+ ua1 = -6.18676573154753e-11 lua1 = 6.32430077202686e-15 wua1 = 9.08755936212857e-15 pua1 = -2.2990715317061e-20
+ ub1 = 4.06081585772902e-19 lub1 = -3.86398114489403e-24 wub1 = -4.98929553461867e-24 pub1 = 1.26308440525738e-29
+ uc1 = -1.20516963553766e-09 luc1 = 4.31503280447514e-15 wuc1 = 7.87239225949609e-15 puc1 = -3.15526689686874e-20
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.12 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.07636237298153 lvth0 = 5.60967311861451e-08 wvth0 = 1.6259851415204e-07 pvth0 = -1.08319576576196e-13
+ k1 = 0.516176246160522 lk1 = -1.80079184353312e-07 wk1 = -6.47106026892919e-07 pk1 = 1.45188329983136e-12
+ k2 = -0.00637185451196262 lk2 = 5.99674128675563e-08 wk2 = 2.22128817622357e-07 pk2 = -4.82161535598342e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 36668.8354567295 lvsat = 0.0334256162433536 wvsat = 0.118214762068338 pvsat = -2.35641977391776e-7
+ ua = -1.2930637317316e-09 lua = 1.41651195929239e-15 wua = 7.44719853142989e-15 pua = -1.88844491489737e-20
+ ub = 1.51150319542223e-18 lub = -8.58238164935004e-25 wub = -4.05045029380802e-24 pub = 9.97218359325022e-30
+ uc = -6.19625728364736e-11 luc = 2.10051914123208e-17 wuc = -1.30919574374239e-16 puc = 4.32201769819667e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00925930203023656 lu0 = 3.72936521545947e-09 wu0 = 2.62887560926926e-08 pu0 = -7.39676062152977e-14
+ a0 = 1.13431230231456 la0 = -3.08491056396393e-07 wa0 = 2.43210953394609e-07 pa0 = 1.55626681645033e-12
+ keta = -0.00909786835714493 lketa = -1.44219659768352e-08 wketa = 2.4935456629057e-08 pketa = -5.38562951121243e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.112013842866754 lags = 1.51490948018711e-06 wags = 1.47075711262695e-06 pags = -5.0506712339144e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.293835593771702 lvoff = 1.12746792244301e-07 wvoff = 3.18688582327384e-08 pvoff = -5.94301130623276e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.33820912601027 lnfactor = 8.05867623585996e-07 wnfactor = 2.26869578289966e-06 pnfactor = -6.90916667143107e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15923519030644 leta0 = -3.16412896387939e-07 weta0 = -3.38841630738418e-14 peta0 = 1.35310916267557e-19
+ etab = -0.139268495046268 letab = 2.76612513471073e-07 wetab = -1.77403851022362e-16 petab = 7.08434150418352e-22
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.02474689264385 lpclm = -2.42707738788853e-06 wpclm = -3.95253957025334e-06 ppclm = 1.62527708408454e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00047479002903789 lpdiblc2 = -7.70693372965986e-10 wpdiblc2 = -3.47783714583786e-09 ppdiblc2 = 1.03734583882938e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 772483502.723579 lpscbe1 = 109.882674200826 wpscbe1 = 197.076679643345 ppscbe1 = -0.000786993793733592
+ pscbe2 = 5.30349045775227e-09 lpscbe2 = 4.66130938903466e-15 wpscbe2 = 2.10686535362533e-14 ppscbe2 = -2.37474838140749e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.949781421168005 lbeta0 = 1.39546182811475e-05 wbeta0 = 2.10212042320702e-05 pbeta0 = -3.90611798923001e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.09958839768263e-10 lagidl = -2.19185133745989e-16 wagidl = -5.55263793440834e-16 pagidl = 1.10682841948977e-21
+ bgidl = -871227871.615888 lbgidl = 2565.8804116806 wbgidl = 12618.291969381 pbgidl = -0.0157990867982182
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.481238919034349 lkt1 = 3.90023030384709e-08 wkt1 = 1.04967608101537e-07 pkt1 = -2.45660865212659e-13
+ kt2 = 0.126050459846816 lkt2 = -3.34261647527979e-07 wkt2 = -9.29574226291119e-07 pkt2 = 1.82113602263992e-12
+ at = 101167.433209994 lat = -0.0330092724137401 wat = 0.0398074474703289 pat = -1.30322123399613e-7
+ ute = -0.326436011397087 lute = 4.82540453957603e-07 wute = 1.05897923393512e-06 pute = -4.22869071285058e-12
+ ua1 = 1.02204857932899e-09 lua1 = 1.99585687541753e-15 wua1 = 9.28594972960573e-15 pua1 = -2.37829551103415e-20
+ ub1 = -3.50091720583559e-19 lub1 = -8.44325546035128e-25 wub1 = -4.7784345592572e-24 pub1 = 1.17888049069457e-29
+ uc1 = 9.61647670837893e-11 luc1 = -8.81635316220402e-16 wuc1 = -2.37392223534164e-15 puc1 = 9.36432806349893e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.06309909752088 lvth0 = 2.96585402059754e-08 wvth0 = 1.19361452997798e-07 pvth0 = -2.21334995691011e-14
+ k1 = 0.327480830921503 lk1 = 1.96054557268403e-07 wk1 = 2.10458031977282e-07 pk1 = -2.57531726148844e-13
+ k2 = 0.0589027282408705 lk2 = -7.01468933678106e-08 wk2 = -4.28998019787076e-08 pk2 = 4.61300829400061e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -72820.2721227911 lvsat = 0.2516744149677 wvsat = 0.765347782150954 pvsat = -1.52559681737722e-6
+ ua = -5.76104297463658e-10 lua = -1.26305254923907e-17 wua = -1.31471736957148e-15 pua = -1.41898923070343e-21
+ ub = 1.06757465867557e-18 lub = 2.66614566465191e-26 wub = 5.85739343906578e-25 pub = 7.30690613187482e-31
+ uc = -5.36881133222912e-11 luc = 4.51139683323947e-18 wuc = 7.63301296754247e-17 puc = 1.90830592487178e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0111350245963138 lu0 = -9.58385295977659e-12 wu0 = -7.36376312989099e-09 pu0 = -6.88676085319117e-15
+ a0 = 0.213430063358942 la0 = 1.52713850403891e-06 wa0 = 7.53860256964215e-06 pa0 = -1.29859145170973e-11
+ keta = -0.0713723724377544 lketa = 1.09712169438199e-07 wketa = 4.53694958222524e-07 pketa = -9.08518902499442e-13
+ a1 = 0.0
+ a2 = 0.44986115912682 la2 = 6.97945056788462e-07 wa2 = 1.76811088061638e-06 pa2 = -3.52444260654609e-12
+ ags = 2.16149251083439 lags = -3.01695712788683e-06 wags = -1.25630468372084e-05 pags = 2.29234434638425e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.22592411111109 lvoff = -2.26237467794384e-08 wvoff = -3.52062325933252e-07 pvoff = 1.71003488159794e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.65671111183595 lnfactor = 1.70985512164207e-07 wnfactor = -2.05207260814041e-06 pnfactor = 1.70358515162794e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.48573896061288 leta0 = 9.69238587657277e-07 weta0 = 6.77683260219522e-14 peta0 = -6.73168551339275e-20
+ etab = 26.0397399007306 letab = -5.190699972415e-05 wetab = -0.000131492735920389 petab = 2.6210946723443e-10
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.49136427670448 lpclm = 2.58838261819793e-06 wpclm = 1.18534330486169e-05 ppclm = -1.52538750073081e-11
+ pdiblc1 = 0.431440277336474 lpdiblc1 = -8.26044795453339e-08 wpdiblc1 = -1.65424453990468e-07 ppdiblc1 = 3.29746850268454e-13
+ pdiblc2 = -0.000251411706063657 lpdiblc2 = 6.7687214127786e-10 wpdiblc2 = 3.44095344768364e-09 ppdiblc2 = -3.41802981581517e-15
+ pdiblcb = -0.0491388386668577 lpdiblcb = 4.81168643905167e-08 wpdiblcb = 3.17788049716879e-10 ppdiblcb = -6.33458995446526e-16
+ drout = 0.646986001581431 ldrout = -1.73392502420327e-07 wdrout = -1.7027703430232e-06 pdrout = 3.39419683002118e-12
+ pscbe1 = 855032994.55284 lpscbe1 = -54.6663647431296 wpscbe1 = -394.153359286687 ppscbe1 = 0.00039152750960712
+ pscbe2 = 2.02894901206716e-09 lpscbe2 = 1.11885772852937e-14 wpscbe2 = 4.8760862227486e-14 ppscbe2 = -7.89474157022394e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000156327218113701 lalpha0 = 3.11613183634129e-10 walpha0 = 7.89412655291583e-10 palpha0 = -1.57356624347361e-15
+ alpha1 = 4.5013884087318e-10 lalpha1 = -6.97945056788463e-16 walpha1 = -1.76811088061638e-15 palpha1 = 3.5244426065461e-21
+ beta0 = -66.4278004856646 lbeta0 = 0.000148260912644149 wbeta0 = 0.000373515344561367 pbeta0 = -7.4170114458802e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -956458108.46995 lbgidl = 2735.7730815508 wbgidl = 12434.6077519975 pbgidl = -0.0154329420677075
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.456094110366761 lkt1 = -1.11197995813612e-08 wkt1 = -2.69716730047349e-09 pkt1 = -3.10485771423662e-14
+ kt2 = -0.036836989935945 lkt2 = -9.57190415291038e-09 wkt2 = -2.56043253981149e-08 pkt2 = 1.92184683336611e-14
+ at = -85625.6790834141 lat = 0.339332536458977 wat = 1.10557266474741 pat = -2.25475243007627e-6
+ ute = 0.292903058864427 lute = -7.52011649679342e-07 wute = -3.24250848702685e-06 pute = 4.3456282178763e-12
+ ua1 = 2.24902479407497e-09 lua1 = -4.49921438531804e-16 wua1 = -5.81802546461183e-15 pua1 = 6.32437259534972e-21
+ ub1 = -4.44619375295072e-19 lub1 = -6.55899979847783e-25 wub1 = 2.92785448511578e-24 pub1 = -3.57243388418665e-30
+ uc1 = -6.77736364354485e-10 luc1 = 6.61011217318505e-16 wuc1 = 4.6267625307692e-15 puc1 = -4.59040290681092e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.02004338370715 lvth0 = -1.31103364423258e-08 wvth0 = -1.2376048801328e-07 pvth0 = 2.19368763070956e-13
+ k1 = 0.5888156193584 lk1 = -6.35392188079261e-08 wk1 = -2.03823373349649e-07 pk1 = 1.53989736455796e-13
+ k2 = -0.0346694007439822 lk2 = 2.2801858093745e-08 wk2 = 1.66456931234654e-08 pk2 = -1.30187200737962e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 184285.666797988 lvsat = -0.00371868418798851 wvsat = -0.98123609241366 pvsat = 2.09351315415046e-7
+ ua = 1.28371693700096e-10 lua = -7.12413297603014e-16 wua = -5.31025976450652e-15 pua = 2.54993486079655e-21
+ ub = 6.4775416056259e-19 lub = 4.4368511060107e-25 wub = 3.20120652400173e-24 pub = -1.86735232455388e-30
+ uc = -8.17040323518775e-11 luc = 3.23406738102506e-17 wuc = 1.68629983503067e-16 puc = -7.2601892952725e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145941945291977 lu0 = -3.44570879575081e-09 wu0 = -2.57790916122185e-08 pu0 = 1.14058847107871e-14
+ a0 = 2.56128558840139 la0 = -8.05075607495703e-07 wa0 = -1.08601880261215e-05 pa0 = 5.29030333571741e-12
+ keta = 0.0783135022673772 lketa = -3.89764979696472e-08 wketa = -8.49566387128427e-07 pketa = 3.8606011576878e-13
+ a1 = 0.0
+ a2 = 1.50658462837287 la2 = -3.51738520705474e-07 wa2 = -3.58068410901885e-06 pa2 = 1.78871871086818e-12
+ ags = -2.44917447063237 lags = 1.5629935901494e-06 wags = 2.00541732918712e-05 pags = -9.47648074473716e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.225907583557786 lvoff = -2.26401642261826e-08 wvoff = -2.39846555175946e-07 pvoff = 5.95352988672683e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.5391686126243 lnfactor = -7.05593056753885e-07 wnfactor = -4.47450545536764e-06 pnfactor = 4.10987975122694e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -52.0813336230975 letab = 2.56936312078623e-05 wetab = 0.00026298492301251 petab = -1.29740181534657e-10
+ dsub = 0.202823170331954 ldsub = 5.67959176287979e-08 wdsub = 1.29387353397984e-07 pdsub = -1.28525374849646e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.60098323812158 lpclm = -4.83363677484353e-07 wpclm = -6.97206050238212e-06 ppclm = 3.4462031056541e-12
+ pdiblc1 = 0.605375734770895 lpdiblc1 = -2.55381178962326e-07 wpdiblc1 = 6.70732757401469e-07 ppdiblc1 = -5.0083988178119e-13
+ pdiblc2 = 0.00043
+ pdiblcb = 0.220612877333715 lpdiblcb = -2.19837765678061e-07 wpdiblcb = -6.35576099433757e-10 ppdiblcb = 3.13553841742194e-16
+ drout = -0.048109443162863 ldrout = 5.17072216471081e-07 wdrout = 3.40554068604641e-06 pdrout = -1.68008263097276e-12
+ pscbe1 = 800000000.0
+ pscbe2 = -2.90988437955433e-09 lpscbe2 = 1.60945081688602e-14 wpscbe2 = 8.20425971828652e-14 ppscbe2 = -1.12007427739346e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000312654736227403 lalpha0 = -1.54244412927155e-10 walpha0 = -1.57882531058317e-09 palpha0 = 7.78894521072479e-16
+ alpha1 = -6.0027768174636e-10 lalpha1 = 3.45473590957386e-16 walpha1 = 3.53622176123277e-15 palpha1 = -1.74455257124305e-21
+ beta0 = 155.296247045962 lbeta0 = -7.19860092828218e-05 wbeta0 = -0.000741516627228073 pbeta0 = 3.65902484205359e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 3074764530.63407 lbgidl = -1268.59355233152 wbgidl = -9730.13787851747 pbgidl = 0.00658414202741697
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.426665543009719 lkt1 = -4.03523138226714e-08 wkt1 = -6.74555518285744e-08 pkt1 = 3.32783870280045e-14
+ kt2 = -0.0378742970358044 lkt2 = -8.54150759295034e-09 wkt2 = -1.24305620973031e-08 pkt2 = 6.13246864395923e-15
+ at = 424290.024863283 lat = -0.167186109068027 wat = -2.24073256849414 pat = 1.06925971770142e-6
+ ute = -0.425714525253207 lute = -3.81814959071009e-08 wute = 1.32530245988015e-06 pute = -1.91751972502409e-13
+ ua1 = 3.09442042783544e-09 lua1 = -1.28968504658016e-15 wua1 = 1.26583890545727e-15 pua1 = -7.12299070285965e-22
+ ub1 = -2.5174169121692e-18 lub1 = 1.40308857983569e-24 wub1 = -1.92863233863185e-24 pub1 = 1.25169902434118e-30
+ uc1 = -4.84160950733e-11 luc1 = 3.58834796712717e-17 wuc1 = 1.10722639565959e-17 puc1 = -5.46236855581912e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.15 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.08819162925908 lvth0 = 2.05097827217694e-08 wvth0 = 6.89351575005131e-07 pvth0 = -1.81770315874422e-13
+ k1 = 0.102010233858814 lk1 = 1.76620376463669e-07 wk1 = 2.36054248865334e-07 pk1 = -6.30186099324991e-14
+ k2 = 0.126991335773725 lk2 = -5.69515263384275e-08 wk2 = -5.51282377039432e-08 pk2 = 2.23900874127359e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 214586.750038586 lvsat = -0.0186673599917385 wvsat = -0.818435157751386 pvsat = 1.29035427910629e-7
+ ua = -5.57954408339692e-10 lua = -3.7382255107491e-16 wua = -5.24481628146432e-16 pua = 1.88928646560936e-22
+ ub = 1.34258818152846e-18 lub = 1.00897084365813e-25 wub = -1.54467818726909e-24 pub = 4.73972947135051e-31
+ uc = -3.19062311658059e-11 luc = 7.77352616871645e-18 wuc = 4.19664632264076e-17 puc = -1.01139651864783e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0112296164664487 lu0 = -1.78583458343032e-09 wu0 = -6.52179043090389e-09 pu0 = 1.90552626059971e-15
+ a0 = 1.2288826280951 la0 = -1.47750595864118e-07 wa0 = -5.01094225701041e-07 pa0 = 1.79768718405565e-13
+ keta = 0.0314663465664558 lketa = -1.58650158704661e-08 wketa = 1.98582715547467e-07 pketa = -1.3103166624714e-13
+ a1 = 0.0
+ a2 = 0.787386106746973 la2 = 3.06943955640516e-09 wa2 = 8.89246955721644e-08 pa2 = -2.16387575711393e-14
+ ags = -0.0476830074917975 lags = 3.78246594706559e-07 wags = -2.04938984343482e-06 pags = 1.42804688530844e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.291202147720405 lvoff = 9.5721254686757e-09 wvoff = 4.99480350440181e-07 pvoff = -3.05202758095579e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.610241922543693 lnfactor = 2.460197786771e-07 wnfactor = 3.48076392060329e-06 pnfactor = 1.85243067824195e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.99636279357148 leta0 = -7.43146007854966e-07 weta0 = -7.26866095849569e-06 peta0 = 3.58590665994235e-12
+ etab = 0.0135140434666189 letab = -6.7367502650702e-09 wetab = -6.16006018278115e-08 petab = 3.06643321931085e-14
+ dsub = 0.233059130242816 ldsub = 4.1879369638293e-08 wdsub = -3.37321844178465e-07 pdsub = 1.01720007264324e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.275271878875414 lpclm = 1.70660113063432e-07 wpclm = 1.42623942752934e-06 ppclm = -6.96997385168564e-13
+ pdiblc1 = -0.371270110801464 lpdiblc1 = 2.26435329200651e-07 wpdiblc1 = 2.60034727413468e-07 ppdiblc1 = -2.98226937062971e-13
+ pdiblc2 = -0.0175397966267037 lpdiblc2 = 8.86518352822473e-09 wpdiblc2 = 6.03900240334085e-08 ppdiblc2 = -2.97926936765937e-14
+ pdiblcb = -0.24812338325364 lpdiblcb = 1.14076436475842e-08 wpdiblcb = -8.66268209748202e-07 ppdiblcb = 4.27363026060758e-13
+ drout = 2.20347302615153 ldrout = -5.93718975775542e-07 wdrout = -4.83921417594755e-06 pdrout = 2.38736824313361e-12
+ pscbe1 = 800012145.528787 lpscbe1 = -0.00599185088026388 wpscbe1 = -0.0613317892493797 ppscbe1 = 3.0257302245304e-8
+ pscbe2 = 6.18965708313068e-08 lpscbe2 = -1.58769788319556e-14 wpscbe2 = -3.70062040175393e-13 ppscbe2 = 1.11032969845702e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.80796803745295e-09 lalpha0 = 3.40796313566097e-15 walpha0 = -6.45731223359516e-15 palpha0 = 3.18563750269736e-21
+ alpha1 = 1.973352e-10 lalpha1 = -4.80191528976e-17
+ beta0 = 3.38890209240018 lbeta0 = 2.95565646187871e-06 wbeta0 = -5.3792309108046e-08 pbeta0 = 1.1069215210608e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -29739831.0699415 lbgidl = 262.976420462822 wbgidl = 3626.32854912971 pbgidl = -5.11040706563382e-6
+ cgidl = 461.556270432166 lcgidl = -7.97018473424639e-05 wcgidl = 0.000466845001557909 pcgidl = -2.30312379378575e-10
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.481728178967838 lkt1 = -1.3187823124365e-08 wkt1 = 1.57660814174172e-07 pkt1 = -7.77800707430581e-14
+ kt2 = 0.0187994330498334 lkt2 = -3.65008122459388e-08 wkt2 = -6.34108329535685e-08 pkt2 = 3.12829735076476e-14
+ at = 17492.6238288657 lat = 0.0335025071634901 wat = 0.323069608566668 pat = -1.95561320725403e-7
+ ute = -0.484655752365456 lute = -9.10354880599812e-09 wute = 7.5678242551706e-07 pute = 8.87205642102133e-14
+ ua1 = 8.99330330902921e-10 lua1 = -2.06763688339668e-16 wua1 = -9.34422304184432e-16 pua1 = 3.73173394356254e-22
+ ub1 = 3.00978003221546e-19 lub1 = 1.26672690666489e-26 wub1 = 9.28744143157988e-25 pub1 = -1.57953374432056e-31
+ uc1 = -4.52399672431535e-11 luc1 = 3.43165751198029e-17 wuc1 = 3.96612237151117e-16 puc1 = -1.95663887851658e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.16 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.71750521473078 lvth0 = -6.96923080167183e-08 wvth0 = -5.17398519924263e-07 pvth0 = 1.11877838725504e-13
+ k1 = 0.42695925292975 lk1 = 9.75479320609852e-08 wk1 = -6.46549873209486e-07 pk1 = 1.51752511924942e-13
+ k2 = 0.0286002974671029 lk2 = -3.30092478589708e-08 wk2 = 2.26240876049351e-07 pk2 = -4.60777099897629e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 310339.438323621 lvsat = -0.0419676276536423 wvsat = -1.07114846853863 pvsat = 1.90530179530974e-7
+ ua = -1.72255887449559e-09 lua = -9.0430029489466e-17 wua = 1.14071420215235e-15 pua = -2.1627677639231e-22
+ ub = 1.40227758887013e-18 lub = 8.63723833621064e-26 wub = -5.62303154072208e-26 pub = 1.11777018891929e-31
+ uc = 1.54233088824656e-13 luc = -2.80030820768359e-20 wuc = -1.43398978647041e-18 puc = 4.47014248769406e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0046405726924412 lu0 = -1.82469849550892e-10 wu0 = 7.55490937453325e-09 pu0 = -1.51986971665575e-15
+ a0 = 0.768832093875613 la0 = -3.58028189682179e-08 wa0 = 1.36304528141361e-06 pa0 = -2.73847260976699e-13
+ keta = -0.220551369452623 lketa = 4.54604711101845e-08 wketa = -4.52696345184815e-08 pketa = -7.16931230867929e-14
+ a1 = 0.0
+ a2 = 0.804864934722957 la2 = -1.18382348561454e-09 wa2 = 4.59669680178922e-07 pa2 = -1.11855100635378e-13
+ ags = 2.14244295756457 lags = -1.54694277378326e-07 wags = 1.32764637083813e-05 pags = -2.30131566628341e-12
+ b0 = 0.0
+ b1 = 1.31755895762121e-23 lb1 = -3.2061216162963e-30 wb1 = -9.28845098453027e-29 pb1 = 2.26023308567363e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.0965116424245087 lvoff = -3.78034727090172e-08 wvoff = -3.71184297167839e-07 pvoff = -9.33369640759381e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.1045437171627 lnfactor = -1.17600631421899e-07 wnfactor = -1.05752118997927e-05 pnfactor = 3.60559611200772e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -3.93148819350829 leta0 = 6.99325395639051e-07 weta0 = 2.47750551522521e-05 peta0 = -4.21154713101481e-12
+ etab = 0.101521044353953 letab = -2.81521978469925e-08 wetab = 1.59902358048617e-07 petab = -2.32357550573018e-14
+ dsub = 0.833221164896261 ldsub = -1.04162859550207e-07 wdsub = -6.04947606141277e-07 pdsub = 1.66843524928832e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.82744607231801 lpclm = -2.07042850820502e-07 wpclm = -5.05802082336134e-06 ppclm = 8.80869535762673e-13
+ pdiblc1 = 1.50803741944381 lpdiblc1 = -2.30871606594175e-07 wpdiblc1 = -3.5394486120025e-06 ppdiblc1 = 6.26331739783834e-13
+ pdiblc2 = 0.0556183270986758 lpdiblc2 = -8.93696798286167e-09 wpdiblc2 = -2.17658331770215e-07 ppdiblc2 = 3.78670371279485e-14
+ pdiblcb = -0.513855059808429 lpdiblcb = 7.60702583570734e-08 wpdiblcb = 3.093815034815e-06 ppdiblcb = -5.36275710504763e-13
+ drout = -3.41358717287403 ldrout = 7.7312521893494e-07 wdrout = 1.89744583258323e-05 pdrout = -3.40740319610449e-12
+ pscbe1 = 799956623.111479 lpscbe1 = 0.00751886310240479 wpscbe1 = 0.219042104465188 ppscbe1 = -3.79683203037551e-8
+ pscbe2 = -3.34073801295645e-08 lpscbe2 = 7.31409398696089e-15 wpscbe2 = 2.92552359326006e-13 ppscbe2 = -5.02062929001691e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.47713144194748e-08 lalpha0 = -4.27647629884293e-15 walpha0 = 2.3061829405697e-14 palpha0 = -3.9974913855247e-21
+ alpha1 = -2.47625714285714e-10 lalpha1 = 6.02567460628571e-17
+ beta0 = 32.5574984252139 lbeta0 = -4.1421714325555e-06 wbeta0 = 2.36719272658651e-06 pbeta0 = -4.78425504509757e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.35193009207452e-11 lagidl = 2.76235596474523e-17 wagidl = 5.73243204373986e-16 pagidl = -1.39491854865957e-22
+ bgidl = 1759526409.76291 lbgidl = -172.420048048964 wbgidl = 8427.5508730041 pbgidl = -0.00117343024491258
+ cgidl = -276.986680114878 lcgidl = 0.000100013717157753 wcgidl = -0.00166730357699253 pcgidl = 2.89007067428731e-10
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.53592367299 wkt1 = -1.619771821234e-7
+ kt2 = -0.131201028226 wkt2 = 6.51468666562244e-8
+ at = 540602.318962161 lat = -0.0937899598308556 wat = -2.34238766058088 pat = 4.53045720234424e-7
+ ute = -1.07196157535862 lute = 1.33810275549513e-07 wute = 3.8982069438669e-06 pute = -6.75707395236002e-13
+ ua1 = -1.60817226263034e-10 lua1 = 5.12104979259819e-17 wua1 = 2.08275628143746e-15 pua1 = -3.61020808311807e-22
+ ub1 = 2.54811740208192e-19 lub1 = 2.39012751757924e-26 wub1 = 9.72076683938877e-25 pub1 = -1.68497828240597e-31
+ uc1 = 9.57843492212001e-11 wuc1 = -4.07470511337231e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.17 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.0161315323171252 lvth0 = -1.91267019378936e-07 wvth0 = -4.89944538177174e-06 pvth0 = 8.71453077664422e-13
+ k1 = -0.392657687757268 lk1 = 2.39618693325791e-07 wk1 = 1.00916539780682e-06 pk1 = -1.35245861722483e-13
+ k2 = 0.803054948003311 lk2 = -1.67251668073616e-07 wk2 = -3.23722795959463e-06 pk2 = 5.54273051043092e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 205485.824211048 lvsat = -0.0237925118905972 wvsat = -0.058712136199623 pvsat = 1.50364905559961e-8
+ ua = -6.21833455280008e-09 lua = 6.88858735036479e-16 wua = 3.7069846718057e-14 pua = -6.44416074843419e-21
+ ub = 4.43901906161463e-18 lub = -4.40010310040481e-25 wub = -2.68906774041579e-23 pub = 4.76320640836179e-30
+ uc = -5.68689044216977e-13 luc = 9.73067946203345e-20 wuc = 5.91137890799853e-18 puc = -8.2621726999245e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0102124660880833 lu0 = 2.39212618658767e-09 wu0 = 1.14522258763292e-07 pu0 = -2.00613761250045e-14
+ a0 = 1.17101362378597 la0 = -1.05516160999819e-07 wa0 = -1.38328229199229e-05 pa0 = 2.36017414130656e-12
+ keta = 0.275607229049946 lketa = -4.05426680370539e-08 wketa = -2.58846860070149e-06 pketa = 3.69139899313439e-13
+ a1 = 0.0
+ a2 = -2.19600370085958 la2 = 5.18980744068992e-07 wa2 = 1.32486678338167e-05 pa2 = -2.32867446259064e-12
+ ags = 1.25
+ b0 = 0.0
+ b1 = -3.07430423444949e-23 lb1 = 4.40664620357521e-30 wb1 = 2.16730522972373e-28 pb1 = -3.1065719701814e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.574511853609982 lvoff = -1.54117343464644e-07 wvoff = -6.80142001570368e-06 pvoff = 1.02126723490363e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -13.723479233335 lnfactor = 2.62599721077148e-06 wnfactor = 9.20303850035655e-05 pnfactor = -1.41798528440266e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.51940007829828 leta0 = 2.81218865924778e-07 weta0 = 6.35996843866777e-06 peta0 = -1.01951283025552e-12
+ etab = -0.231132122977319 letab = 2.95092368718757e-08 wetab = -1.11565828990309e-07 petab = 2.38199975476516e-14
+ dsub = 0.0999383576860371 ldsub = 2.29429156859987e-08 wdsub = 2.06610389251714e-06 pdsub = -2.96151199745622e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.71862137087371 lpclm = -5.3485539472155e-07 wpclm = -1.12835390361757e-05 ppclm = 1.95998841173549e-12
+ pdiblc1 = 0.924450429477843 lpdiblc1 = -1.29713804927454e-07 wpdiblc1 = 4.27021779990339e-07 ppdiblc1 = -6.12083050234236e-14
+ pdiblc2 = 0.0339848896858175 lpdiblc2 = -5.18707120859164e-09 wpdiblc2 = -8.40619177647916e-08 ppdiblc2 = 1.47097019170764e-14
+ pdiblcb = -1.28618179332612 lpdiblcb = 2.09943829691563e-07 wpdiblcb = 6.11615581363059e-06 ppdiblcb = -1.0601622164231e-12
+ drout = 1.26942818544336 ldrout = -3.861929724508e-08 wdrout = -3.94695129404574e-06 pdrout = 5.65748104585929e-13
+ pscbe1 = 1037237333.48986 lpscbe1 = -41.1222449124662 wpscbe1 = -1197.98737433922 ppscbe1 = 0.000207656735493214
+ pscbe2 = 1.14644682539838e-08 lpscbe2 = -4.63902468146611e-16 wpscbe2 = -9.38564160314656e-15 ppscbe2 = 2.13103630488838e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 18.6713885325858 lbeta0 = -1.73518091598713e-06 wbeta0 = -2.95954589535218e-05 pbeta0 = 5.06191661241687e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.37890482199508e-10 lagidl = -1.19958109339046e-16 wagidl = -4.67218093371007e-15 pagidl = 7.69739474381258e-22
+ bgidl = -1130940033.82741 lbgidl = 328.607624350096 wbgidl = 13478.3817633864 pbgidl = -0.00204893116978967
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.164051748335465 lkt1 = -1.21332339581714e-07 wkt1 = -6.8075615838838e-07 pkt1 = 8.9924110187821e-14
+ kt2 = -0.175354045021279 lkt2 = 7.65339562526016e-09 wkt2 = 3.76414252415214e-07 pkt2 = -5.39544661126921e-14
+ at = -184329.302219754 lat = 0.0318682375215751 wat = 1.56736426415516 pat = -2.24662858895472e-7
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.71945786510145e-10 luc1 = -4.78692712167912e-17 wuc1 = -2.35433744980576e-15 puc1 = 3.37466021380258e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.18 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0537489431687 wvth0 = 5.86524686695862e-8
+ k1 = 0.44205207135451 wk1 = -5.80141215968923e-8
+ k2 = 0.0248237253676165 wk2 = -5.31710770688974e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 323282.33637695 wvsat = -0.822955660079779
+ ua = -1.10744223691828e-09 wua = 2.78940299102583e-15
+ ub = 1.2393304653032e-18 wub = -8.11355992844838e-25
+ uc = -9.27767945288183e-12 wuc = -2.72434533704855e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00853738103508001 wu0 = 1.26067771702569e-8
+ a0 = 1.3101985775754 wa0 = -5.83783413380071e-7
+ keta = -0.012282397655245 wketa = 3.7473305957607e-8
+ a1 = 0.0
+ a2 = 1.07716489714687 wa2 = -8.45281483187463e-7
+ ags = 0.309122196092176 wags = -4.08481756909438e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.278390185468769 wvoff = -5.73912519381443e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.41438576175584 wnfactor = 1.51744570432627e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.347005573953947 wpclm = -6.04564498173483e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000133338415931977 wpdiblc2 = 1.78567236809097e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 865373846.835292 wpscbe1 = -330.121073140511
+ pscbe2 = 7.8629967022153e-09 wpscbe2 = 6.13072686726336e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.25320264185616e-10 walpha0 = -6.32835026573253e-16
+ alpha1 = 2.5248701384693e-10 walpha1 = -7.70020108774829e-16
+ beta0 = 1.27556883885757 wbeta0 = 2.56304465703625e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1831914799.42999 wbgidl = -1461.96803056708
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.423448049072474 wkt1 = -6.36549844626647e-8
+ kt2 = -0.0472892886219128 wkt2 = -1.63933688432524e-8
+ at = 90000.0
+ ute = -0.154755494649972 wute = -5.0278340702204e-8
+ ua1 = 1.72985419276207e-09 wua1 = 1.15892950575362e-15
+ ub1 = -7.7370399143252e-19 wub1 = 1.07442513567083e-25
+ uc1 = 1.1396316068919e-10 wuc1 = -1.02636045017316e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.19 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0537489431687 wvth0 = 5.86524686695879e-8
+ k1 = 0.44205207135451 wk1 = -5.80141215968931e-8
+ k2 = 0.0248237253676165 wk2 = -5.3171077068898e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 323282.33637695 wvsat = -0.822955660079779
+ ua = -1.10744223691828e-09 wua = 2.78940299102583e-15
+ ub = 1.2393304653032e-18 wub = -8.11355992844838e-25
+ uc = -9.2776794528818e-12 wuc = -2.72434533704855e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00853738103508001 wu0 = 1.26067771702568e-8
+ a0 = 1.3101985775754 wa0 = -5.83783413380071e-7
+ keta = -0.012282397655245 wketa = 3.7473305957607e-8
+ a1 = 0.0
+ a2 = 1.07716489714687 wa2 = -8.45281483187465e-7
+ ags = 0.309122196092176 wags = -4.08481756909438e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.278390185468769 wvoff = -5.73912519381438e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.41438576175584 wnfactor = 1.51744570432627e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.347005573953947 wpclm = -6.04564498173483e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000133338415931977 wpdiblc2 = 1.78567236809097e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 865373846.835292 wpscbe1 = -330.12107314051
+ pscbe2 = 7.8629967022153e-09 wpscbe2 = 6.13072686726336e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.25320264185616e-10 walpha0 = -6.32835026573253e-16
+ alpha1 = 2.5248701384693e-10 walpha1 = -7.70020108774829e-16
+ beta0 = 1.27556883885757 wbeta0 = 2.56304465703625e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1831914799.42999 wbgidl = -1461.96803056707
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.423448049072474 wkt1 = -6.36549844626656e-8
+ kt2 = -0.0472892886219128 wkt2 = -1.63933688432524e-8
+ at = 90000.0
+ ute = -0.154755494649972 wute = -5.02783407022042e-8
+ ua1 = 1.72985419276207e-09 wua1 = 1.15892950575362e-15
+ ub1 = -7.7370399143252e-19 wub1 = 1.07442513567083e-25
+ uc1 = 1.1396316068919e-10 wuc1 = -1.02636045017318e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.20 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.06262269978816 lvth0 = 7.09309359890674e-08 wvth0 = 6.99529191074277e-08 pvth0 = -9.03283199018835e-14
+ k1 = 0.530793050435021 lk1 = -7.09336640241456e-07 wk1 = -4.27339440244663e-07 pk1 = 2.95214210390933e-12
+ k2 = -0.00610486988431966 lk2 = 2.47222715713921e-07 wk2 = 1.25899871399314e-07 pk2 = -1.04886166533482e-12
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 548343.001603383 lvsat = -1.79898596765972 wvsat = -1.43743032144168 pvsat = 4.91170366070124e-6
+ ua = -1.64119992627694e-09 lua = 4.26650562114275e-15 wua = 4.70334052511315e-15 pua = -1.52987496208464e-20
+ ub = 1.44675049405168e-18 lub = -1.65797839775631e-24 wub = -1.40676265850699e-24 pub = 4.75928672609059e-30
+ uc = 5.95594457962296e-12 luc = -1.21767505856734e-16 wuc = -3.59605785576392e-16 puc = 6.96789280092326e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00587205428747613 lu0 = 2.13048575740384e-08 wu0 = 2.25511735555569e-08 pu0 = -7.94889215136818e-14
+ a0 = 1.32862577376842 la0 = -1.47294807563097e-07 wa0 = -6.15368556722904e-07 pa0 = 2.52470726517685e-13
+ keta = -0.0129741666777652 lketa = 5.52954361493362e-09 wketa = 6.91001360601783e-08 pketa = -2.52803942878427e-13
+ a1 = 0.0
+ a2 = 1.35386817615754 la2 = -2.21178283484059e-06 wa2 = -1.68915515006468e-06 pa2 = 6.74536744864898e-12
+ ags = 0.348472695282173 lags = -3.14541840494371e-07 wags = -1.0100218765759e-06 pags = 4.8083134970545e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.277638024913813 lvoff = -6.01227354603256e-09 wvoff = -6.61957634316593e-08 pvoff = 7.03774362925567e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.4504189948289 lnfactor = -2.8802581118571e-07 wnfactor = 1.67945572669866e-06 pnfactor = -1.29500086821006e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.212075360148291 lpclm = 1.07854280536088e-06 wpclm = -9.96685515937816e-07 ppclm = 3.13435583189431e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000322784426404387 lpdiblc2 = -1.51430599445751e-09 wpdiblc2 = -4.69556414514648e-10 ppdiblc2 = 5.18067141082484e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 930638813.52868 lpscbe1 = -521.684938338991 wpscbe1 = -659.692329633705 ppscbe1 = 0.00263437444823481
+ pscbe2 = 6.3331713917849e-09 lpscbe2 = 1.22284107872252e-14 wpscbe2 = 1.18984913767618e-14 ppscbe2 = -4.61036912288251e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.20364460368239e-10 lalpha0 = 3.96134149739854e-17 walpha0 = -6.07809494901723e-16 palpha0 = -2.00037533280245e-22
+ alpha1 = 2.53834796508647e-10 lalpha1 = -1.0773282365639e-17 walpha1 = -7.76826063758127e-16 palpha1 = 5.44022985942843e-23
+ beta0 = -9.69692649132035 lbeta0 = 8.77068638775337e-05 wbeta0 = 7.94311761784672e-05 pbeta0 = -4.30047416404189e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.54406130953349e-10 lagidl = -4.34886593982381e-16 wagidl = -2.74736935413853e-16 pagidl = 2.1960651858471e-21
+ bgidl = 1435802806.08597 lbgidl = 3166.25704865253 wbgidl = 819.438396469894 pbgidl = -0.0182360526866788
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.368870747285083 lkt1 = -4.36254820314618e-07 wkt1 = -2.04077764051027e-07 pkt1 = 1.12244674014928e-12
+ kt2 = -0.0431578686030913 lkt2 = -3.30238366304066e-08 wkt2 = -3.27594345306962e-08 pkt2 = 1.30819494769942e-13
+ at = 12613.5593365334 lat = 0.618575976840033 wat = 0.368994300011135 pat = -2.9494961600624e-6
+ ute = -0.027887934724782 lute = -1.0140952877173e-06 wute = -4.84842005339567e-07 pute = 3.47361425396509e-12
+ ua1 = 1.27911773946639e-09 lua1 = 3.60288882011355e-15 wua1 = 2.31592881441541e-15 pua1 = -9.24828653990001e-21
+ ub1 = -6.24466392744989e-19 lub1 = -1.19290656861779e-24 wub1 = 2.14706081627819e-25 pub1 = -8.57393954595471e-31
+ uc1 = 3.57861121649557e-10 luc1 = -1.94955883946702e-15 wuc1 = -2.05101149701663e-17 puc1 = 8.19038214947304e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.21 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.05461346271302 lvth0 = 3.89473452259103e-08 wvth0 = 5.27721241651509e-08 pvth0 = -2.17195985887146e-14
+ k1 = 0.373015378371156 lk1 = -7.92770668372826e-08 wk1 = 7.58194485716647e-08 pk1 = 9.42858593161316e-13
+ k2 = 0.0458286860643386 lk2 = 3.98344732690177e-08 wk2 = -4.14704549886032e-08 pk2 = -3.8049538089755e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 98301.1165003386 lvsat = -0.00181660628610292 wvsat = -0.193012368399835 pvsat = -5.76778390629876e-8
+ ua = 1.15223286153522e-10 lua = -2.74748593713789e-15 wua = 3.35712147503249e-16 pua = 2.14266674934153e-21
+ ub = 6.77593851070971e-19 lub = 1.41352405261099e-24 wub = 1.60576913336901e-25 pub = -1.49962994505735e-30
+ uc = -6.04314185481519e-11 luc = 1.43339674041208e-16 wuc = -1.38651508798689e-16 puc = -1.85555829626594e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0143527239856468 lu0 = -1.25613229971153e-08 wu0 = 5.68288302050885e-10 pu0 = 8.29616951878358e-15
+ a0 = 1.03422763702158 la0 = 1.02833645903724e-06 wa0 = 7.48612711297419e-07 pa0 = -5.19436750235606e-12
+ keta = -0.0141123846217396 lketa = 1.00748325828883e-08 wketa = 5.02574710229668e-08 pketa = -1.77558812564059e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.332223406673803 lags = -2.496529388216e-07 wags = -7.72526473189937e-07 pags = 3.85991407788799e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.275784622900298 lvoff = -1.34135342358804e-08 wvoff = -5.92838911275679e-08 pvoff = 4.27759939694741e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.63005129719678 lnfactor = -1.00535831025887e-06 wnfactor = 7.94968055319523e-07 pnfactor = 2.23705736043976e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.280058625165649 leta0 = -7.98901710101742e-07 weta0 = -6.1012723164166e-07 peta0 = 2.43644425894945e-12
+ etab = -0.244894021371516 letab = 6.98410941515688e-07 wetab = 5.33381677504415e-07 petab = -2.12997332128213e-12
+ dsub = 1.31493822630977 ldsub = -3.0147235067754e-06 wdsub = -2.30236696717005e-06 pdsub = 9.19412949994492e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0135958562374929 lpclm = 1.97972424926045e-06 wpclm = 1.29082362683677e-06 ppclm = -6.00044135329489e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000867982236533001 lpdiblc2 = 3.24082776978356e-09 wpdiblc2 = 3.30281662860508e-09 ppdiblc2 = -9.88368921244079e-15
+ pdiblcb = 0.0109618223819394 lpdiblcb = -1.43607711867049e-07 wpdiblcb = -1.81597932070984e-07 ppdiblcb = 7.2518192286048e-13
+ drout = 0.56
+ pscbe1 = 829062731.07521 lpscbe1 = -116.057308386416 wpscbe1 = -88.6338374073166 ppscbe1 = 0.000353944871004461
+ pscbe2 = 8.69514328830249e-09 lpscbe2 = 2.79625865792938e-15 wpscbe2 = 3.94168111007434e-15 ppscbe2 = -1.4329458432072e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.84803028897529e-10 lalpha0 = -2.17711569399633e-16 walpha0 = -9.33207653711671e-16 palpha0 = 1.09938729942555e-21
+ alpha1 = 4.01770528127303e-10 lalpha1 = -6.01530660996222e-16 walpha1 = -1.52386337060073e-15 palpha1 = 3.03757476342652e-21
+ beta0 = 13.6788228296188 lbeta0 = -5.64040416424703e-06 wbeta0 = -4.32571733337314e-05 pbeta0 = 5.9888631860156e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.07229865515796e-11 lagidl = -1.40644893483307e-16 wagidl = 9.73439483004568e-17 pagidl = 7.10220453837163e-22
+ bgidl = 2584536810.133 lbgidl = -1421.02610160067 wbgidl = -4832.42877731601 pbgidl = 0.00433376326935304
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.505091761503496 lkt1 = 1.07721732162309e-07 wkt1 = 2.25418313307938e-07 pkt1 = -5.92676266419217e-13
+ kt2 = -0.0753600598698912 lkt2 = 9.55703974385738e-08 wkt2 = 8.74969746462684e-08 pkt2 = -3.4940499373998e-13
+ at = 175682.251731657 lat = -0.0326124291117261 wat = -0.336473176143857 pat = -1.32326079768581e-7
+ ute = -1.41237058533168 lute = 4.51461189129194e-06 wute = 6.54266887837163e-06 pute = -2.45896120033724e-11
+ ua1 = 3.14777222840417e-10 lua1 = 7.4538264500957e-15 wua1 = 1.28574877453173e-14 pua1 = -5.13442943979099e-20
+ ub1 = 4.71851051745124e-19 lub1 = -5.57087267976306e-24 wub1 = -8.92903366267034e-24 pub1 = 3.56566494284207e-29
+ uc1 = -5.31956518410092e-10 luc1 = 1.6037837556535e-15 wuc1 = 7.97928326735067e-16 puc1 = -3.18639750842756e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.22 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.02932531166733 lvth0 = -1.14604872032017e-08 wvth0 = -5.11874586806516e-08 pvth0 = 1.85506988361975e-13
+ k1 = 0.10039887683441 lk1 = 4.6413976510297e-07 wk1 = 1.35716335838934e-06 pk1 = -1.61129291334682e-12
+ k2 = 0.162272482600208 lk2 = -1.92277371230199e-07 wk2 = -5.64890412770687e-07 pk2 = 6.62857510907873e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 244068.671580339 lvsat = -0.292380612994161 wvsat = -0.834859689580168 pvsat = 1.22174081644397e-6
+ ua = -1.73563971923514e-09 lua = 9.41909624297528e-16 wua = 4.54063758214276e-15 pua = -6.2391709066919e-21
+ ub = 1.62637248106967e-18 lub = -4.77712444153367e-25 wub = -2.23604560110502e-24 pub = 3.27764878463528e-30
+ uc = 5.31004707896902e-11 luc = -8.2967755187707e-17 wuc = -4.62924689993097e-16 puc = 4.60830224829106e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00595722128274793 lu0 = 4.17375156967585e-09 wu0 = 1.87828087659224e-08 pu0 = -2.80115262736291e-14
+ a0 = 3.05232777324131 la0 = -2.99441923029471e-06 wa0 = -6.79709899743419e-06 pa0 = 9.84678638370358e-12
+ keta = 0.10088003799562 lketa = -2.19143933132354e-07 wketa = -4.16135307794606e-07 pketa = 7.52119636378603e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = -1.64763899562792 lags = 3.69688202245772e-06 wags = 6.67208527632395e-06 pags = -1.09797134176645e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.313009896080735 lvoff = 6.07890173550665e-08 wvoff = 8.76984374480882e-08 pvoff = -2.50209466908865e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.214745534570712 lnfactor = 1.81582444800265e-06 wnfactor = 5.22948181832324e-06 pnfactor = -6.60242743487854e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.727385830331298 leta0 = 1.20927560592963e-06 weta0 = 1.22025446328332e-06 peta0 = -1.21212512804893e-12
+ etab = -34.2820315755331 letab = 6.8545930639453e-05 wetab = 0.000173116659082056 petab = -3.46146778336317e-10
+ dsub = -0.65187505261954 ldsub = 9.0580014101899e-07 wdsub = 4.60473393434011e-06 pdsub = -4.57405719686954e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.8471449765229 lpclm = -1.72936116083248e-06 wpclm = -5.0051780124959e-06 ppclm = 6.54961796244923e-12
+ pdiblc1 = 0.390866386212638 lpdiblc1 = -1.72700056032672e-09 wpdiblc1 = 3.94632362357761e-08 ppdiblc1 = -7.86635683917507e-14
+ pdiblc2 = 0.00108351045437734 lpdiblc2 = -6.49156767730276e-10 wpdiblc2 = -3.30005931961042e-09 ppdiblc2 = 3.27807432442317e-15
+ pdiblcb = -0.121021474460452 lpdiblcb = 1.19479609094169e-07 wpdiblcb = 3.6330656746386e-07 ppdiblcb = -3.60996922433307e-13
+ drout = 0.230293343769541 ldrout = 6.57216806717111e-07 wdrout = 4.01420155559661e-07 pdrout = -8.00166050042983e-13
+ pscbe1 = 741874537.849581 lpscbe1 = 57.7382303215727 wpscbe1 = 177.267674814635 ppscbe1 = -0.00017608671756502
+ pscbe2 = 1.32054628524648e-08 lpscbe2 = -6.19433272145884e-15 wpscbe2 = -7.67765136125417e-15 ppscbe2 = 8.83179851766105e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.5066333061691e-10 lalpha0 = -1.4965961150834e-16 walpha0 = -7.6081097860876e-16 palpha0 = 7.55742455869269e-22
+ alpha1 = 1.0e-10
+ beta0 = 12.673999595604 lbeta0 = -3.63745182860242e-06 wbeta0 = -2.59283534049786e-05 pbeta0 = 2.53464366010158e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.90704969165552e-11 lagidl = 1.77877529266097e-16 wagidl = 9.04259845054499e-16 pagidl = -8.98235665966746e-22
+ bgidl = 2578052665.42636 lbgidl = -1408.10100955941 wbgidl = -5413.76045930138 pbgidl = 0.00549255380165839
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391249452887838 lkt1 = -1.19204467609008e-07 wkt1 = -3.30145970616336e-07 pkt1 = 5.14751132169828e-13
+ kt2 = -0.0110141705813727 lkt2 = -3.26927088240231e-08 wkt2 = -1.56002906015875e-07 pkt2 = 1.35972571379336e-13
+ at = 351979.590328345 lat = -0.384032613435371 wat = -1.10422113114352 pat = 1.39805509335454e-6
+ ute = 1.6847753734155 lute = -1.65904683982524e-06 wute = -1.02711048508271e-05 pute = 8.92592209444106e-12
+ ua1 = 3.686021553228e-09 lua1 = 7.33797019049587e-16 wua1 = -1.30744886405701e-14 pua1 = 3.46899547182051e-22
+ ub1 = -7.5076055188382e-19 lub1 = -3.13379451100854e-24 wub1 = 4.47378850369363e-24 pub1 = 8.94029469696506e-30
+ uc1 = 7.14555127546979e-10 luc1 = -8.80935275675275e-16 wuc1 = -2.40395057058658e-15 puc1 = 3.19602936900178e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.08326102983466 lvth0 = 4.21159112097006e-08 wvth0 = 1.95472327421469e-07 pvth0 = -5.9509550245132e-14
+ k1 = 0.606367207056303 lk1 = -3.84578041029854e-08 wk1 = -2.92454366424754e-07 pk1 = 2.73350581845565e-14
+ k2 = -0.0564653548022676 lk2 = 2.50032346995016e-08 wk2 = 1.26709642120851e-07 pk2 = -2.41351044179779e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -131455.051406357 lvsat = 0.080641370949998 wvsat = 0.613173136561131 pvsat = -2.16645215009572e-7
+ ua = -1.85246834309527e-11 lua = -7.63765991138129e-16 wua = -4.56847092988074e-15 pua = 2.80925272442449e-21
+ ub = 8.33963468675203e-19 lub = 3.0941753940053e-25 wub = 2.26089752279267e-24 pub = -1.189335704171e-30
+ uc = -4.1567900070096e-11 luc = 1.10699349854114e-17 wuc = -3.40471374250269e-17 puc = 3.48098545162443e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0138438141188205 lu0 = -3.66030078492281e-09 wu0 = -2.19898639878834e-08 pu0 = 1.24895189342909e-14
+ a0 = -0.66051158659657 la0 = 6.93685193727924e-07 wa0 = 5.40905712830643e-06 pa0 = -2.27805232992735e-12
+ keta = -0.221735743270409 lketa = 1.01322581798881e-07 wketa = 6.65604950141895e-07 pketa = -3.22414067959525e-13
+ a1 = 0.0
+ a2 = 0.855668795604156 la2 = -5.52979300878407e-08 wa2 = -2.93726959638508e-07 pa2 = 2.91770150633396e-13
+ ags = 3.4206042760025 lags = -1.33759661249711e-06 wags = -9.58669614967402e-06 pags = 5.17075200647346e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.27415565940833 lvoff = 2.21936276073727e-08 wvoff = 3.79378951534595e-09 pvoff = -1.66863791740651e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.2574641838547 lnfactor = -2.13285609639805e-07 wnfactor = -3.0519707134829e-06 pnfactor = 1.62385406016071e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 68.9839487907733 letab = -3.40320917656531e-05 wetab = -0.000348363542547731 petab = 1.71859322190214e-10
+ dsub = 0.224453312887367 ldsub = 3.53098750830884e-08 wdsub = 2.01607097438947e-08 pdsub = -2.00263990955808e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.406119044464942 lpclm = 5.08891615247537e-07 wpclm = 3.16328859371136e-06 ppclm = -1.56443031922749e-12
+ pdiblc1 = 1.00904408541858 lpdiblc1 = -6.15786399934154e-07 wpdiblc1 = -1.36768834766852e-06 ppdiblc1 = 1.31911357166057e-12
+ pdiblc2 = 0.000666837698516518 lpdiblc2 = -2.35259885769001e-10 wpdiblc2 = -1.19596932074974e-09 ppdiblc2 = 1.1880017731349e-15
+ pdiblcb = 0.220530859393146 lpdiblcb = -2.19797303111296e-07 wpdiblcb = -2.21406643782003e-10 ppdiblcb = 1.09228310830117e-16
+ drout = 0.785275872460918 ldrout = 1.05931571631876e-07 wdrout = -8.02840311119321e-07 pdrout = 3.96071633406984e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 2.53824092974694e-08 lpscbe2 = -1.82901563492468e-14 wpscbe2 = -6.0826192132795e-14 ppscbe2 = 6.16262637105818e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.57425481733679 lbeta0 = 4.3498044995201e-07 wbeta0 = -6.08391403110394e-07 pbeta0 = 1.95156186004012e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.6182827825113e-10 lagidl = -1.60750178261421e-16 wagidl = -8.17191085838074e-16 pagidl = 8.11746958824222e-22
+ bgidl = 772337411.716175 lbgidl = 385.584569130557 wbgidl = 1896.52550630667 pbgidl = -0.00176903103884678
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.514009554323414 lkt1 = 2.73780603080502e-09 wkt1 = 3.73609188019475e-07 pkt1 = -1.84315609599152e-13
+ kt2 = -0.0328143309139654 lkt2 = -1.10377811595661e-08 wkt2 = -3.79820865533236e-08 pkt2 = 1.87380066160436e-14
+ at = -134217.756003195 lat = 0.0989256861749088 wat = 0.579587741575663 pat = -2.7453624465459e-7
+ ute = 0.342407017985139 lute = -3.25621342378752e-07 wute = -2.55351331173964e-06 pute = 1.25974515018701e-12
+ ua1 = 8.51884992919061e-09 lua1 = -4.06683505427237e-15 wua1 = -2.61261316584609e-14 pua1 = 1.33115925192877e-20
+ ub1 = -8.24516964542902e-18 lub1 = 4.31068682915546e-24 wub1 = 2.69950423496756e-23 pub1 = -1.3430922555895e-29
+ uc1 = -3.66276989096027e-10 luc1 = 1.92696337406656e-16 wuc1 = 1.61618783423289e-15 puc1 = -7.97326873764784e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.951832437393914 lvth0 = -2.27228077278341e-08 wvth0 = 7.7280948571156e-10 pvth0 = 3.65431205342582e-14
+ k1 = 0.163421034192796 lk1 = 1.80064374925152e-07 wk1 = -7.40544611169513e-08 pk1 = -8.04099143001847e-14
+ k2 = 0.113533628240646 lk2 = -5.88637235969233e-08 wk2 = 1.28297159411033e-08 pk2 = 3.20461906036865e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 25456.3242167981 lvsat = 0.00323102672282168 wvsat = 0.136624734824863 pvsat = 1.84542204061952e-8
+ ua = -9.29658715624296e-10 lua = -3.1426894996393e-16 wua = 1.3525292982704e-15 pua = -1.11801686131143e-22
+ ub = 1.02857980744732e-18 lub = 2.13405904063373e-25 wub = 4.09831504818267e-26 pub = -9.41675875639128e-32
+ uc = -4.75896127117167e-11 luc = 1.40406746566033e-17 wuc = 1.21163496857495e-16 puc = -4.17614493794266e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00899873800679532 lu0 = -1.27004062596853e-09 wu0 = 4.74357066987863e-09 pu0 = -6.99100252900136e-16
+ a0 = 0.571238059801894 la0 = 8.60162866729989e-08 wa0 = 2.81984130340993e-06 pa0 = -1.00069377330456e-12
+ keta = 0.101631076408027 lketa = -5.8206558287639e-08 wketa = -1.55731081685113e-07 pketa = 8.27822073099479e-14
+ a1 = 0.0
+ a2 = 0.688662408791688 la2 = 2.70926667694481e-08 wa2 = 5.87453919277015e-07 pa2 = -1.4294986180903e-13
+ ags = -2.81930579041722 lags = 1.74078813985027e-06 wags = 1.19465906859851e-05 pags = -5.45243665445695e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.0860307542340639 lvoff = -7.06155368614891e-08 wvoff = -5.36582293480602e-07 pvoff = 9.97242642924044e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.58868573574939 lnfactor = 1.16648212391568e-07 wnfactor = -1.46012509327047e-06 pnfactor = 8.38536125576345e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.366482927314561 leta0 = 6.09356656044893e-08 weta0 = 9.61812183072228e-07 peta0 = -4.74498498772486e-13
+ etab = 0.00464865828736444 letab = -1.98179689275993e-09 wetab = -1.68326921688757e-08 petab = 6.65304348992104e-15
+ dsub = 0.294072112845111 ldsub = 9.6427554953515e-10 wdsub = -6.45421677173141e-07 pdsub = 3.08330684501296e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.794166853835649 lpclm = -8.32550292482797e-08 wpclm = -1.19404642489531e-06 ppclm = 5.85208624181893e-13
+ pdiblc1 = -0.801818314507566 lpdiblc1 = 2.77580834720609e-07 wpdiblc1 = 2.43419216080237e-06 ppdiblc1 = -5.56498554627437e-13
+ pdiblc2 = -0.0043274684194413 lpdiblc2 = 2.22862110585207e-09 wpdiblc2 = -6.32882727505457e-09 ppdiblc2 = 3.72023565059574e-15
+ pdiblcb = -0.567731063497013 lpdiblcb = 1.6908225740349e-07 wpdiblcb = 7.47668180620868e-07 ppdiblcb = -3.68853124891138e-13
+ drout = 1.00440263087424 ldrout = -2.17198511023697e-09 wdrout = 1.21578219985483e-06 pdrout = -5.99791558911982e-13
+ pscbe1 = 800000000.0
+ pscbe2 = -4.3110488492554e-08 lpscbe2 = 1.54999928606878e-14 wpscbe2 = 1.60196538590211e-13 ppscbe2 = -4.74126482188446e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.05703849742862e-08 lalpha0 = 1.01974863824444e-14 walpha0 = 6.30393453463266e-14 palpha0 = -3.10997045544661e-20
+ alpha1 = 3.4575883349272e-10 lalpha1 = -1.21242171397631e-16 walpha1 = -7.49501085525521e-16 palpha1 = 3.6975736653099e-22
+ beta0 = -6.47112278601071 lbeta0 = 7.85743694603227e-06 wbeta0 = 4.97367914124534e-05 pbeta0 = -2.46420356138606e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.43185516096839e-09 lagidl = -1.72464490052739e-15 wagidl = -1.68250096106299e-14 pagidl = 8.70901213420795e-21
+ bgidl = 213203934.577475 lbgidl = 661.42636047521 wbgidl = 2399.52516351304 pbgidl = -0.00201717988373366
+ cgidl = 586.270015136891 lcgidl = -0.000141227876727604 wcgidl = -0.000162927257997569 pcgidl = 8.03782076060047e-11
+ egidl = 1.97886865382484 legidl = -9.26917303940642e-07 wegidl = -9.48780232947651e-06 pegidl = 4.68069342561929e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.400324591436112 lkt1 = -5.33473061900915e-08 wkt1 = -2.53406317016177e-07 pkt1 = 1.25014965624127e-13
+ kt2 = 0.0915056319202278 lkt2 = -7.23695429842614e-08 wkt2 = -4.30558393590991e-07 pkt2 = 2.12410816777392e-13
+ at = 66816.0075095094 lat = -0.000251908648921745 wat = 0.0739992365477296 pat = -2.51102227611195e-8
+ ute = -0.33479019576 lute = 8.46577665584692e-9
+ ua1 = 4.29498206488999e-10 lua1 = -7.60504540981951e-17 wua1 = 1.4381088013842e-15 pua1 = -2.86894740691394e-22
+ ub1 = 5.51281263333473e-19 lub1 = -2.89366692716141e-26 wub1 = -3.35222792226797e-25 pub1 = 5.21357886808695e-32
+ uc1 = 1.17907496082509e-11 luc1 = 6.18115532976476e-18 wuc1 = 1.08621819570329e-16 puc1 = -5.35872712231869e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.25 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.872075470773442 lvth0 = -4.21307084713266e-08 wvth0 = 2.63141424879187e-07 pvth0 = -2.73011335983598e-14
+ k1 = 0.5872654990847 lk1 = 7.69269105272855e-08 wk1 = -1.45605508934173e-06 pk1 = 2.55883354570775e-13
+ k2 = -0.0286485264068586 lk2 = -2.42654024493088e-08 wk2 = 5.15332677866063e-07 pk2 = -9.02318751452093e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -56002.2210168059 lvsat = 0.0230529862028764 wvsat = 0.778782468250751 pvsat = -1.37807158130194e-7
+ ua = -1.94484830035453e-09 lua = -6.72347467948452e-17 wua = 2.26321849652601e-15 pua = -3.3340697425626e-22
+ ub = 1.74686672431862e-18 lub = 3.8619402285744e-26 wub = -1.79631661434303e-24 pub = 3.52917262609037e-31
+ uc = 3.47284410300679e-11 luc = -5.99043590481514e-18 wuc = -1.76024826658942e-16 puc = 3.05557628884162e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00513970925320032 lu0 = -3.30992287126226e-10 wu0 = 5.034398420105e-09 pu0 = -7.69869695984721e-16
+ a0 = 3.33141756518768 la0 = -5.85640273808568e-07 wa0 = -1.15773507141778e-05 pa0 = 2.50269013787121e-12
+ keta = -0.0806582499923219 lketa = -1.3848638180031e-08 wketa = -7.51693823346802e-07 pketa = 2.2780258894042e-13
+ a1 = 0.0
+ a2 = 0.558328548562314 la2 = 5.88078476499434e-08 wa2 = 1.7046148732098e-06 pa2 = -4.14797574017127e-13
+ ags = 11.9724486774532 lags = -1.85860780885238e-06 wags = -3.63625310015815e-05 pags = 6.30300839875213e-12
+ b0 = 0.0
+ b1 = -1.31755895762121e-23 lb1 = 3.2061216162963e-30 wb1 = 4.01821515404542e-29 pb1 = -9.77784439155104e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.0961063178566346 lvoff = -6.81637693607001e-08 wvoff = -3.73231081742935e-07 pvoff = 5.99747071305837e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -2.06280383418596 lnfactor = 1.0051943813605e-06 wnfactor = 1.04688188923193e-05 pnfactor = -2.06422924598909e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.59573856023088 leta0 = -2.38188941598102e-07 weta0 = -3.13601503507358e-06 peta0 = 5.22658580836678e-13
+ etab = 0.0406813692995357 letab = -1.07499247250397e-08 wetab = 4.67127032605198e-07 petab = -1.11112748017153e-13
+ dsub = 0.166883633834733 ldsub = 3.19140656549622e-08 wdsub = 2.75988514390392e-06 pdsub = -5.20309866725955e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0335155624375654 lpclm = 1.18151554562812e-07 wpclm = 4.33935567624487e-06 ppclm = -7.61278376305355e-13
+ pdiblc1 = 0.66815501043113 lpdiblc1 = -8.01195342233238e-08 wpdiblc1 = 7.01741031826505e-07 ppdiblc1 = -1.34927361804708e-13
+ pdiblc2 = 0.00562324910435547 lpdiblc2 = -1.92766594953582e-10 wpdiblc2 = 3.48039233699959e-08 ppdiblc2 = -6.28892562586955e-15
+ pdiblcb = 0.910068479288695 lpdiblcb = -1.90522527738899e-07 wpdiblcb = -4.0966317501371e-06 ppdiblcb = 8.09949131659644e-13
+ drout = 1.53850669319406 ldrout = -1.32139799427018e-07 wdrout = -6.03233904801292e-06 pdrout = 1.16395176930166e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 4.8803272583498e-08 lpscbe2 = -6.86611793203657e-15 wpscbe2 = -1.2259024296869e-13 ppscbe2 = 2.14001216321354e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.39228034795937e-08 lalpha0 = -1.27962971095458e-14 walpha0 = -2.25140519094024e-13 palpha0 = 3.90254072987199e-20
+ alpha1 = -7.77710119616857e-10 lalpha1 = 1.52140516714147e-16 walpha1 = 2.67678959116258e-15 palpha1 = -4.63989354152939e-22
+ beta0 = 68.4900003161139 lbeta0 = -1.03834528273925e-05 wbeta0 = -0.000179082678423471 pbeta0 = 3.10384365370736e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.21942749144563e-08 lagidl = 2.0777863397663e-15 wagidl = 6.20829188539313e-14 pagidl = -1.04922853625014e-20
+ bgidl = 7131481718.19918 lbgidl = -1022.05351883573 wbgidl = -18699.4385445206 pbgidl = 0.00311699974705182
+ cgidl = -722.392911203183 lcgidl = 0.000177219542442137 wcgidl = 0.000581883064277032 pcgidl = -1.00862446595652e-10
+ egidl = -6.61024519223159 legidl = 1.16314048113104e-06 wegidl = 3.3885008319559e-05 pegidl = -5.87355957209572e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.860500726041802 lkt1 = 5.86310340525878e-08 wkt1 = 1.47705325982393e-06 pkt1 = -2.96071606884989e-13
+ kt2 = -0.436632348495648 lkt2 = 5.6146496894177e-08 wkt2 = 1.60749629382358e-06 pkt2 = -2.83525334748695e-13
+ at = 153765.342308894 lat = -0.0214099858803345 wat = -0.38896065505447 pat = 8.75455113415765e-8
+ ute = -0.3
+ ua1 = 7.32574130346422e-11 lua1 = 1.06364680994012e-17 wua1 = 9.00739697426206e-16 pua1 = -1.56132417672464e-22
+ ub1 = 5.30588259791808e-19 lub1 = -2.39012751757925e-26 wub1 = -4.20523644771641e-25 pub1 = 7.28927275374267e-32
+ uc1 = 3.7192270660305e-11 wuc1 = -1.11595619642564e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.26 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.58932328220464 lvth0 = 8.21955926665348e-08 wvth0 = 3.04476738632712e-06 pvth0 = -5.09462614503821e-13
+ k1 = -0.0350215001207808 lk1 = 1.84792894395565e-07 wk1 = -7.96805151148258e-07 pk1 = 1.41610288784197e-13
+ k2 = -0.159538280445407 lk2 = -1.57723426377513e-09 wk2 = 1.62361968753711e-06 pk2 = -2.82340128827568e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169619.735154785 lvsat = -0.0160558724359948 wvsat = 0.122402367256745 pvsat = -2.40315441840944e-8
+ ua = 6.45831239663715e-09 lua = -1.52382181568999e-15 wua = -2.69439523370175e-14 pua = 4.7293056036885e-21
+ ub = -5.18513091974681e-18 lub = 1.24019800991276e-24 wub = 2.17087988958522e-23 pub = -3.72141244969719e-30
+ uc = 7.31852179223179e-13 luc = -9.7535186587409e-20 wuc = -6.56018990846856e-19 puc = 1.576845048439e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0285603820110996 lu0 = -4.39068486163497e-09 wu0 = -8.12706284973415e-08 pu0 = 1.41900710598316e-14
+ a0 = -5.61744441828076 la0 = 9.65537564681884e-07 wa0 = 2.04471401280309e-05 pa0 = -3.04837105573556e-12
+ keta = -0.705107081218503 lketa = 9.43920733270528e-08 wketa = 2.36388583800499e-06 pketa = -3.12245758398976e-13
+ a1 = 0.0
+ a2 = 2.44215683986062 la2 = -2.67731180707122e-07 wa2 = -1.01728471790329e-05 pa2 = 1.64401794319453e-12
+ ags = 1.25
+ b0 = 0.0
+ b1 = 3.07430423444949e-23 lb1 = -4.40664620357521e-30 wb1 = -9.3758353594393e-29 pb1 = 1.34391348875131e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.980044083558183 lvoff = 8.50562350704748e-08 wvoff = 1.04868670247494e-06 pvoff = -1.86497677750175e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 15.3361089942057 lnfactor = -2.01069837048726e-06 wnfactor = -5.47130439836701e-05 pnfactor = 9.23426450120916e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.149907636831496 leta0 = 1.24284990021005e-08 weta0 = -2.06960517520864e-06 peta0 = 3.37809228547409e-13
+ etab = -0.0502303205623976 letab = 5.00852577224816e-09 wetab = -1.025073294701e-06 petab = 1.47542272317449e-13
+ dsub = 0.785782032553578 ldsub = -7.53645449821647e-08 wdsub = -1.39722985506456e-06 pdsub = 2.00276132965244e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.41917561129315 lpclm = -1.33655028109323e-07 wpclm = 3.28069252589311e-07 ppclm = -6.59700102017489e-14
+ pdiblc1 = 1.09673359026096 lpdiblc1 = -1.54408488093867e-07 wpdiblc1 = -4.42963767365563e-07 ppdiblc1 = 6.34934786776462e-14
+ pdiblc2 = 0.0114313462497088 lpdiblc2 = -1.19953053793484e-09 wpdiblc2 = 2.98276622840598e-08 ppdiblc2 = -5.42635048175556e-15
+ pdiblcb = -0.188015344889178 lpdiblcb = -1.82873823554952e-10 wpdiblcb = 5.70698356334438e-07 ppdiblcb = 9.23465664080792e-16
+ drout = -0.293204208071499 ldrout = 1.85365304776552e-07 wdrout = 3.94393944657323e-06 pdrout = -5.65316392392914e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.03975245252142e-08 lpscbe2 = -2.08942375109786e-16 wpscbe2 = -3.99785083095377e-15 ppscbe2 = 8.43553563764412e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.5299447529672 lbeta0 = -3.36772716187804e-07 wbeta0 = 1.15167332693456e-05 pbeta0 = -1.99968428693587e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.98817400935598e-10 lagidl = 1.19854325287652e-16 wagidl = 4.09774615282994e-15 pagidl = -4.41251496837919e-22
+ bgidl = 2358841974.44934 lbgidl = -194.773690933619 wbgidl = -4144.11771260946 pbgidl = 0.000594009544690016
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.278988308483013 lkt1 = -1.38885716213875e-07 wkt1 = -1.26115615648829e-06 pkt1 = 1.78564136919738e-13
+ kt2 = -0.0685659549787205 lkt2 = -7.65339562526016e-09 wkt2 = -1.62838072330096e-07 pkt2 = 2.33408836116513e-14
+ at = -6781.76583984483 lat = 0.00641892875195169 wat = 0.670794977191492 pat = -9.61504104406741e-8
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.34046627238648e-11 luc1 = 6.56536384486661e-19 wuc1 = -6.44792050586758e-16 puc1 = 9.24232029470047e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.034517
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29720858
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.911951
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.28 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.034517
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29720858
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.911951
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.29 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0396853777065 lvth0 = 4.13125899197166e-8
+ k1 = 0.390669914700905 lk1 = 2.58660623235218e-7
+ k2 = 0.0351772658317135 lk2 = -9.66954244275052e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77014.5327768425 lvsat = -0.188455195353381
+ ua = -9.89907109822351e-11 lua = -7.49901870889343e-16
+ ub = 9.85477846643321e-19 lub = -9.74246151806612e-26
+ uc = -1.11957558265434e-10 luc = 1.06707307552848e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0132665066958 lu0 = -4.75928696699256e-9
+ a0 = 1.126848536098 la0 = -6.45105228725166e-8
+ keta = 0.00968353076963815 lketa = -7.73640015766657e-08 wketa = -2.99852972050473e-24 pketa = 4.18096279767136e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.017289988568175 lags = 1.26208765200978e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.299343388544765 lvoff = 1.70642462635953e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.00110676335525 lnfactor = -7.12652151146524e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.114734399685775 lpclm = 2.10628732484659e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168818489705 lpdiblc2 = 1.84418379958414e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714327962.84966 lpscbe1 = 342.117401489868
+ pscbe2 = 1.02346458760091e-08 lpscbe2 = -2.88883132878883e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1065813124638e-11 lalpha0 = -2.59782056161896e-17
+ alpha1 = -8.83803561262884e-13 lalpha1 = 7.06504462287938e-18 walpha1 = 2.34440593327997e-34 palpha1 = -2.72457263015603e-39
+ beta0 = 16.3482835524884 lbeta0 = -5.33042079449267e-05 wbeta0 = 1.35525271560688e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.43208327881951e-11 lagidl = 2.85195643082475e-16
+ bgidl = 1704493843.79725 lbgidl = -2813.28203720162
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435787145678045 lkt1 = -6.82083867015476e-8
+ kt2 = -0.0538995747481865 lkt2 = 9.87142670363557e-9
+ at = 133605.523841315 lat = -0.348553690730689
+ ute = -0.18686596419218 lute = 1.24890903956571e-7
+ ua1 = 2.0385028489407e-09 lua1 = 5.70407405815647e-16
+ ub1 = -5.54065005497301e-19 lub1 = -1.47404310356671e-24
+ uc1 = 3.51135925346025e-10 luc1 = -1.92270285751067e-15 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.30 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0373096643247 lvth0 = 3.1825563395068e-8
+ k1 = 0.39787631532893 lk1 = 2.29883029764101e-7
+ k2 = 0.0322306662092167 lk2 = -8.4928656184203e-08 pk2 = 5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35013.023362553 lvsat = -0.0207289717519407
+ ua = 2.2530214708257e-10 lua = -2.04491286412814e-15
+ ub = 7.3024646981917e-19 lub = 9.21800540683538e-25
+ uc = -1.05894772401041e-10 luc = 8.24965543747024e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145390637694 lu0 = -9.84103748616824e-9
+ a0 = 1.279695175654 la0 = -6.74878816783792e-7
+ keta = 0.00236686763209579 lketa = -4.81460926363186e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0789146275940702 lags = 1.01599963925139e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29522360732579 lvoff = 6.12567370175419e-10
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.8907185940324 lnfactor = -2.71834879839156e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.40966078061423 lpclm = 1.22001243377312e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0485835162604495 lpdiblcb = 9.41769516564709e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.9876069955871e-09 lpscbe2 = -1.90232158012222e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.1192557782444e-11 lalpha0 = 1.42773752745155e-16
+ alpha1 = -9.78990408614235e-11 lalpha1 = 3.94479678312628e-16 walpha1 = -2.00296714216273e-32 palpha1 = 5.87747175411144e-38
+ beta0 = -0.5050558384638 lbeta0 = 1.39968726718593e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1264173309365e-10 lagidl = 9.223395569849e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43117787025461 lkt1 = -8.66147814024163e-8
+ kt2 = -0.046670102192069 lkt2 = -1.89983007746655e-8
+ at = 65353.85212337 lat = -0.0760016964958941
+ ute = 0.73294808402065 lute = -3.54823748770556e-06 pute = 8.07793566946316e-28
+ ua1 = 4.5307033248294e-09 lua1 = -9.38179145816879e-15
+ ub1 = -2.45594843985464e-18 lub1 = 6.12082028642297e-24
+ uc1 = -2.7031855873761e-10 luc1 = 5.5897494905091e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.31 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0461095036822 lvth0 = 4.93666175802695e-8
+ k1 = 0.5454080839698 lk1 = -6.41976508749532e-8
+ k2 = -0.0229531449202714 lk2 = 2.50713315250285e-08 wk2 = -2.64697796016969e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -29678.9552125639 lvsat = 0.108224007437026
+ ua = -2.46780240508461e-10 lua = -1.10389310181221e-15
+ ub = 8.93180803063241e-19 lub = 5.97017342723469e-25
+ uc = -9.86909462006041e-11 luc = 6.81368938639756e-17 wuc = 9.86076131526265e-32
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0121160398104 lu0 = -5.01113175378311e-9
+ a0 = 0.823582341108001 la0 = 2.34308228604462e-7
+ keta = -0.0355693011631478 lketa = 2.74735141976547e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.540114866427681 lags = 9.6671677575281e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.28425387944166 lvoff = -2.12538080709204e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.9294746740774 lnfactor = -3.49088846923895e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32726858 leta0 = 8.1182393672004e-07 peta0 = -2.01948391736579e-28
+ etab = 22.482326763364 letab = -4.49544099258305e-05 wetab = 6.67038445962762e-21 petab = 1.81753552562921e-26
+ dsub = 0.858001400000001 ldsub = -5.940175146732e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.20596428508744 lpclm = 4.18236089338113e-7
+ pdiblc1 = 0.40380624592792 lpdiblc1 = -2.75205146454682e-8
+ pdiblc2 = 1.43233000000041e-06 lpdiblc2 = 4.2571255218246e-10
+ pdiblcb = -0.00189449793638372 lpdiblcb = 1.10995724841425e-9
+ drout = 0.361917635016081 ldrout = 3.94845105252317e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.06879873224826e-08 lpscbe2 = -3.29841630017542e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.19602200021408e-12 lalpha0 = 9.81457458983515e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.17218150587221 lbeta0 = 4.67355773837533e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.1743320265992e-10 lagidl = -1.166508626638e-16
+ bgidl = 802899192.027401 lbgidl = 392.888530362486
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499503183520001 lkt1 = 4.95806618913891e-8
+ kt2 = -0.0621669880280001 lkt2 = 1.18922306437575e-8
+ at = -10090.7286459999 lat = 0.0743848532457603
+ ute = -1.6830846545 lute = 1.26773237923172e-06 pute = 1.61558713389263e-27
+ ua1 = -6.0105839752e-10 lua1 = 8.47544189935722e-16 wua1 = 3.94430452610506e-31
+ ub1 = 7.16179343460001e-19 lub1 = -2.02302564913869e-25
+ uc1 = -7.3692013666e-11 luc1 = 1.67031784950957e-16 wuc1 = 2.46519032881566e-32 puc1 = -4.70197740328915e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.32 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0191663245768 lvth0 = 2.26029339340693e-8
+ k1 = 0.510472424072761 lk1 = -2.94947323441472e-8
+ k2 = -0.014917698045952 lk2 = 1.70894167977859e-08 wk2 = 6.61744490042422e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 69602.315528176 lvsat = 0.0096041485219607
+ ua = -1.5165106213508e-09 lua = 1.57378335232961e-16
+ ub = 1.5753040065058e-18 lub = -8.05615559377584e-26
+ uc = -5.27318395745652e-11 luc = 2.24839668062795e-17 puc = 2.35098870164458e-38
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0066334131912 lu0 = 4.34969606879774e-10
+ a0 = 1.113099680712 la0 = -5.32803464830964e-8
+ keta = -0.00348616462015639 lketa = -4.39588448968728e-9
+ a1 = 0.0
+ a2 = 0.75935673367364 la2 = 4.03725008860937e-8
+ ags = 0.27715951215524 lags = 3.57875223277559e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.27291168884736 lvoff = -3.25204369914811e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.2567334619324 lnfactor = 3.19170563265793e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.243261151015 letab = 2.2319990121863e-5
+ dsub = 0.23106394041644 ldsub = 2.87432875546143e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.63111242831704 lpclm = -4.07971696129197e-9
+ pdiblc1 = 0.5605837704226 lpdiblc1 = -1.83253587271965e-7
+ pdiblc2 = 0.00027468346307008 lpdiblc2 = 1.54281818160893e-10
+ pdiblcb = 0.220458260914565 lpdiblcb = -2.1976148752307e-07 wpdiblcb = -1.65436122510606e-23 ppdiblcb = -2.60324098722934e-29
+ drout = 0.52202728996784 ldrout = 2.35802100821846e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.43770966587601e-09 lpscbe2 = 1.91688400668287e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3747653643888 lbeta0 = 4.98971493524154e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.12587401724004e-12 lagidl = 1.05418863444537e-16
+ bgidl = 1394201615.9452 lbgidl = -194.474636807173
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.39150438388 lkt1 = -5.76986497454087e-8
+ kt2 = -0.045268526732 lkt2 = -4.89365310308857e-9
+ at = 55827.075188 lat = 0.00890619382090246
+ ute = -0.494881232720001 lute = 8.74447686476191e-8
+ ua1 = -4.78189710399998e-11 lua1 = 2.97990444514932e-16
+ ub1 = 6.0641208816e-19 lub1 = -9.32665790686782e-26
+ uc1 = 1.6366545464e-10 luc1 = -6.87444079011883e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.33 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.951579035816 lvth0 = -1.07404439286061e-8
+ k1 = 0.1391388305636 lk1 = 1.53698240010475e-7
+ k2 = 0.117740448063352 lk2 = -4.8355887687486e-08 pk2 = 1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70255.10584 lvsat = 0.00928210225510609
+ ua = -4.861690008968e-10 lua = -3.50928339118574e-16
+ ub = 1.0420180418272e-18 lub = 1.82528675304853e-25
+ uc = -7.860517951676e-12 luc = 3.47238739486535e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01055413854848 lu0 = -1.49927319943003e-9
+ a0 = 1.49585434488 la0 = -2.42107766994409e-7
+ keta = 0.050567389226496 lketa = -3.10625566372871e-08 pketa = 6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.88128653265272 la2 = -1.97801022826473e-8
+ ags = 1.097940292214 lags = -4.70471251950703e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.26197424659896 lvoff = -3.79162928754222e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.1099157291336 lnfactor = 3.91601329929288e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.68185784099488 leta0 = -9.4650763560732e-8
+ etab = -0.000870723701341264 letab = 1.99713232889716e-10
+ dsub = 0.0824405601279197 ldsub = 1.02064848739392e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.402643129340079 lpclm = 1.08632870057404e-7
+ pdiblc1 = -0.00365505965856028 lpdiblc1 = 9.51068686826147e-8
+ pdiblc2 = -0.00640266916101696 lpdiblc2 = 3.44847360702274e-09 wpdiblc2 = -8.27180612553028e-25 ppdiblc2 = -1.18329135783152e-30
+ pdiblcb = -0.3225732332316 lpdiblcb = 4.8136583736011e-8
+ drout = 1.40305344137712 ldrout = -1.98841578662106e-07 wdrout = -1.6940658945086e-21
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4174066817368e-09 lpscbe2 = -4.64517597278701e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.8374004106232 lbeta0 = -2.22601954915029e-07 wbeta0 = 1.35525271560688e-20
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.08500774325672e-09 lagidl = 1.1310102870514e-15 pagidl = 1.88079096131566e-37
+ bgidl = 1000000000.0
+ cgidl = 532.846726441352 lcgidl = -0.000114872138329124
+ egidl = -1.1321491658048 legidl = 6.07866005159808e-07 wegidl = 4.2351647362715e-22
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.48341565304 lkt1 = -1.23553280405526e-8
+ kt2 = -0.049672987568 lkt2 = -2.72076520317801e-9
+ at = 91080.103192 lat = -0.00848546450853489 wat = 1.11022302462516e-16
+ ute = -0.33479019576 lute = 8.46577665584692e-9
+ ua1 = 9.01049146559999e-10 lua1 = -1.70122254885617e-16 wua1 = -7.88860905221012e-31 pua1 = -1.88079096131566e-37
+ ub1 = 4.4136286032e-19 lub1 = -1.18415231045482e-26
+ uc1 = 4.74074714316e-11 luc1 = -1.13899269811227e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.34 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.785792300714286 lvth0 = -5.10826564747872e-8
+ k1 = 0.109830032788 lk1 = 1.60830184243594e-7
+ k2 = 0.140327289931343 lk2 = -5.38521246139591e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 199357.877371429 lvsat = -0.0221335079638087
+ ua = -1.20274672320286e-09 lua = -1.76557749328064e-16
+ ub = 1.15786067182571e-18 lub = 1.54339761406275e-25
+ uc = -2.29894954758249e-11 luc = 4.02869387225787e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679047121599999 lu0 = -5.83429918079006e-10
+ a0 = -0.464755998 la0 = 2.34983232621324e-7
+ keta = -0.327136074690686 lketa = 6.08470488653921e-8
+ a1 = 0.0
+ a2 = 1.117265914878 la2 = -7.72028531945827e-8
+ ags = 0.0492995661671429 lags = 2.0812701179972e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.218487508549715 lvoff = -4.84982687388495e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.36988594933714 lnfactor = 3.28340696485398e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.567449993717428 leta0 = -6.68109868199316e-8
+ etab = 0.193850720008982 letab = -4.71834134366929e-08 wetab = 5.02512222125964e-23 petab = 7.34626717987067e-30
+ dsub = 1.07184049999343 ldsub = -1.38693753827601e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.38934427018857 lpclm = -1.31469012154387e-7
+ pdiblc1 = 0.898253486238858 lpdiblc1 = -1.24361753058971e-7
+ pdiblc2 = 0.0170353361227257 lpdiblc2 = -2.25488372271263e-9
+ pdiblcb = -0.433203011048126 lpdiblcb = 7.50570126103288e-8
+ drout = -0.439476576346856 ldrout = 2.49515990790811e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.60635267050002e-09 lpscbe2 = 1.50908501258472e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.76940471184571 lbeta0 = -2.06056017565912e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.16250109563771e-09 lagidl = -1.36259801878749e-15
+ bgidl = 1000000000.0
+ cgidl = -531.595451576257 lcgidl = 0.000144147092385325 wcgidl = -2.16840434497101e-19 pcgidl = -2.58493941422821e-26
+ egidl = 4.50053273501714 legidl = -7.62779543222401e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.376180031714286 lkt1 = -3.84498296627092e-8
+ kt2 = 0.0904601689714285 lkt2 = -3.68204872491695e-8
+ at = 26226.4785142858 lat = 0.00729588681329076
+ ute = -0.3
+ ua1 = 3.68606868285714e-10 lua1 = -4.05588157749091e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.35 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = 0.563947705288165 lvth0 = -2.85043889635241e-07 wvth0 = -3.52215401226537e-06 pvth0 = 6.10523132178055e-13
+ k1 = 1.1621400030665 lk1 = -2.15751213845409e-08 wk1 = -4.44783910763394e-06 pk1 = 7.70979535239053e-13
+ k2 = 0.196801235004252 lk2 = -6.3641205305007e-08 wk2 = 5.36876029742731e-07 pk2 = -9.30610172435454e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 166575.3705211 lvsat = -0.0164510537913863 wvsat = 0.131686894552284 pvsat = -2.28263429279037e-8
+ ua = -9.19908293852142e-09 lua = 1.20951117756283e-15 wua = 2.08070669586988e-14 pua = -3.60665537248692e-21
+ ub = 6.49203981318285e-18 lub = -7.70276182598288e-25 wub = -1.39035614649683e-23 pub = 2.41001553721467e-30
+ uc = -3.94304914786051e-13 luc = 1.12088730788524e-19 wuc = 2.77846982258246e-18 puc = -4.81614402106797e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0202401630908956 lu0 = 4.10200617140966e-09 wu0 = 6.75584532832165e-08 pu0 = -1.17104471752062e-14
+ a0 = -1.65176677274049 la0 = 4.40737306293291e-07 wa0 = 8.35284566083008e-06 pa0 = -1.44786556115696e-12
+ keta = -0.450576214903672 lketa = 8.22439158896306e-08 wketa = 1.58763231380209e-06 pketa = -2.75197010009826e-13
+ a1 = 0.0
+ a2 = -0.893484834715332 la2 = 2.71336660238426e-7
+ ags = -10.3645163606705 lags = 2.0132370369259e-06 wags = 3.54212806777271e-05 pags = -6.13985395011586e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.296966117646507 lvoff = -1.3784596939645e-07 wvoff = -2.84586519796949e-06 pvoff = 4.93296581685636e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -16.1671722290247 lnfactor = 3.36817928700628e-06 wnfactor = 4.13638422012832e-05 pnfactor = -7.16992567948602e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.01574925099338 leta0 = 2.0761760385975e-07 weta0 = 1.48534782631153e-06 peta0 = -2.57467221517188e-13
+ etab = -0.250295517592581 letab = 2.98040070966869e-08 wetab = -4.14926020566733e-07 petab = 7.19224465529963e-14
+ dsub = 0.330562837006492 ldsub = -1.02021662807714e-08 wdsub = -8.92866415455878e-09 pdsub = 1.54767678722307e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.43122109036495 lpclm = -3.12065856410121e-07 wpclm = -2.75840855325518e-06 ppclm = 4.78137021804147e-13
+ pdiblc1 = 0.95148729129 lpdiblc1 = -1.33589194358926e-7
+ pdiblc2 = 0.0212117343376133 lpdiblc2 = -2.97881223648482e-9
+ pdiblcb = -0.245247273470374 lpdiblcb = 4.24771409700764e-08 wpdiblcb = 7.45240984115895e-07 ppdiblcb = -1.29178581704681e-13
+ drout = 1.0
+ pscbe1 = 617872337.420839 lpscbe1 = 31.5696447761463 wpscbe1 = 555.442418355022 ppscbe1 = -9.62792779128233e-5
+ pscbe2 = 6.53942374298324e-09 lpscbe2 = 5.09185827696371e-16 wpscbe2 = 7.76836193646916e-15 ppscbe2 = -1.34655232134369e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 14.9251119737245 lbeta0 = -1.09973600292546e-06 wbeta0 = -1.88739367985472e-06 pbeta0 = 3.27157045678659e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.68430126385546e-10 lagidl = 1.85471737375578e-16 wagidl = 3.70009857929166e-15 pagidl = -6.41367687537257e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.279092992818759 lkt1 = -5.5278702810782e-08 wkt1 = 4.40847939122636e-07 pkt1 = -7.64157000716393e-14
+ kt2 = -0.102764678099045 lkt2 = -3.3272787076678e-09 wkt2 = -5.85407832439275e-08 pkt2 = 1.01473422859359e-14
+ at = 94560.1438756112 lat = -0.00454893407311069 wat = 0.361728278503676 pat = -6.27012563392702e-8
+ ute = 0.55761956064625 lute = -1.486580594033e-07 wute = -2.61551856564833e-06 pute = 4.5336875713235e-13
+ ua1 = 1.39125024527775e-10 lua1 = -7.80891941595511e-19 wua1 = -1.37391634143906e-17 pua1 = 2.38151910792368e-24
+ ub1 = 3.04264409813457e-19 lub1 = 1.53292483317552e-26 wub1 = 2.69705751373809e-25 pub1 = -4.67502555316328e-32
+ uc1 = -4.86875125689353e-10 luc1 = 8.4498041338841e-17 wuc1 = 9.41927175944102e-16 puc1 = -1.63271772823799e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.36 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.034517
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29720858
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.911951
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.034517
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29720858
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.911951
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.38 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0396853777065 lvth0 = 4.13125899197166e-8
+ k1 = 0.390669914700905 lk1 = 2.58660623235217e-7
+ k2 = 0.0351772658317135 lk2 = -9.66954244275053e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77014.5327768425 lvsat = -0.18845519535338
+ ua = -9.89907109822347e-11 lua = -7.49901870889345e-16
+ ub = 9.8547784664332e-19 lub = -9.74246151806642e-26
+ uc = -1.11957558265435e-10 luc = 1.06707307552848e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0132665066958 lu0 = -4.75928696699256e-9
+ a0 = 1.126848536098 la0 = -6.45105228725098e-8
+ keta = 0.00968353076963815 lketa = -7.73640015766658e-08 wketa = -5.98413474393831e-24 pketa = 3.44140569902666e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0172899885681752 lags = 1.26208765200978e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.299343388544765 lvoff = 1.70642462635944e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.00110676335525 lnfactor = -7.12652151146537e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.114734399685775 lpclm = 2.1062873248466e-06 ppclm = 1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168818489705 lpdiblc2 = 1.84418379958414e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714327962.849661 lpscbe1 = 342.117401489864
+ pscbe2 = 1.02346458760091e-08 lpscbe2 = -2.88883132878889e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1065813124638e-11 lalpha0 = -2.59782056161897e-17 walpha0 = 4.93038065763132e-32
+ alpha1 = -8.83803561262885e-13 lalpha1 = 7.06504462287938e-18 walpha1 = -5.98843842082906e-34 palpha1 = -5.57183174346062e-39
+ beta0 = 16.3482835524884 lbeta0 = -5.33042079449269e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.43208327881949e-11 lagidl = 2.85195643082476e-16
+ bgidl = 1704493843.79725 lbgidl = -2813.28203720161
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435787145678044 lkt1 = -6.82083867015476e-8
+ kt2 = -0.0538995747481865 lkt2 = 9.87142670363578e-9
+ at = 133605.523841315 lat = -0.348553690730689
+ ute = -0.18686596419218 lute = 1.2489090395657e-7
+ ua1 = 2.0385028489407e-09 lua1 = 5.70407405815647e-16
+ ub1 = -5.54065005497301e-19 lub1 = -1.4740431035667e-24
+ uc1 = 3.51135925346025e-10 luc1 = -1.92270285751067e-15 wuc1 = 3.94430452610506e-31
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.39 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0373096643247 lvth0 = 3.18255633950646e-8
+ k1 = 0.397876315328929 lk1 = 2.29883029764102e-7
+ k2 = 0.0322306662092167 lk2 = -8.49286561842029e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35013.0233625529 lvsat = -0.0207289717519407
+ ua = 2.25302147082569e-10 lua = -2.04491286412813e-15 pua = -1.50463276905253e-36
+ ub = 7.30246469819168e-19 lub = 9.21800540683538e-25
+ uc = -1.05894772401041e-10 luc = 8.24965543747022e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145390637694 lu0 = -9.84103748616821e-9
+ a0 = 1.279695175654 la0 = -6.74878816783794e-7
+ keta = 0.00236686763209581 lketa = -4.81460926363185e-08 pketa = 5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0789146275940702 lags = 1.01599963925139e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29522360732579 lvoff = 6.12567370176266e-10
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.8907185940324 lnfactor = -2.71834879839156e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.40966078061423 lpclm = 1.22001243377312e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0485835162604495 lpdiblcb = 9.41769516564709e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.98760699558709e-09 lpscbe2 = -1.90232158012223e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.1192557782444e-11 lalpha0 = 1.42773752745155e-16 palpha0 = -9.4039548065783e-38
+ alpha1 = -9.78990408614235e-11 lalpha1 = 3.94479678312628e-16 walpha1 = 4.00593428432545e-32 palpha1 = 3.58525777000798e-37
+ beta0 = -0.505055838463804 lbeta0 = 1.39968726718594e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1264173309365e-10 lagidl = 9.2233955698489e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431177870254609 lkt1 = -8.66147814024155e-8
+ kt2 = -0.046670102192069 lkt2 = -1.89983007746655e-8
+ at = 65353.85212337 lat = -0.0760016964958941
+ ute = 0.73294808402065 lute = -3.54823748770555e-06 wute = -4.2351647362715e-22 pute = 8.07793566946316e-28
+ ua1 = 4.5307033248294e-09 lua1 = -9.38179145816879e-15
+ ub1 = -2.45594843985464e-18 lub1 = 6.12082028642296e-24
+ uc1 = -2.7031855873761e-10 luc1 = 5.5897494905091e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.40 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0461095036822 lvth0 = 4.93666175802686e-8
+ k1 = 0.5454080839698 lk1 = -6.41976508749527e-8
+ k2 = -0.0229531449202714 lk2 = 2.50713315250286e-08 wk2 = 2.64697796016969e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -29678.9552125641 lvsat = 0.108224007437026
+ ua = -2.46780240508459e-10 lua = -1.10389310181221e-15
+ ub = 8.93180803063238e-19 lub = 5.97017342723469e-25
+ uc = -9.8690946200604e-11 luc = 6.81368938639755e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0121160398104 lu0 = -5.01113175378311e-9
+ a0 = 0.823582341107999 la0 = 2.34308228604462e-7
+ keta = -0.0355693011631478 lketa = 2.74735141976547e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.540114866427679 lags = 9.66716775752801e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.28425387944166 lvoff = -2.12538080709206e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.9294746740774 lnfactor = -3.49088846923894e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32726858 leta0 = 8.1182393672004e-07 peta0 = 4.03896783473158e-28
+ etab = 22.482326763364 letab = -4.49544099258305e-05 wetab = -1.52465930505774e-20 petab = 1.85792520397653e-26
+ dsub = 0.8580014 ldsub = -5.94017514673199e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.20596428508744 lpclm = 4.18236089338114e-7
+ pdiblc1 = 0.40380624592792 lpdiblc1 = -2.75205146454677e-8
+ pdiblc2 = 1.43232999999954e-06 lpdiblc2 = 4.2571255218246e-10
+ pdiblcb = -0.00189449793638372 lpdiblcb = 1.10995724841425e-09 wpdiblcb = -3.30872245021211e-24
+ drout = 0.36191763501608 ldrout = 3.94845105252317e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.06879873224826e-08 lpscbe2 = -3.29841630017542e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.19602200021382e-12 lalpha0 = 9.81457458983515e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.1721815058722 lbeta0 = 4.67355773837533e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.1743320265992e-10 lagidl = -1.16650862663799e-16
+ bgidl = 802899192.027399 lbgidl = 392.888530362485
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499503183519999 lkt1 = 4.95806618913891e-8
+ kt2 = -0.0621669880279999 lkt2 = 1.18922306437576e-8
+ at = -10090.728646 lat = 0.0743848532457603
+ ute = -1.6830846545 lute = 1.26773237923172e-6
+ ua1 = -6.0105839752e-10 lua1 = 8.47544189935722e-16 wua1 = -7.88860905221012e-31 pua1 = -7.52316384526264e-37
+ ub1 = 7.16179343459999e-19 lub1 = -2.0230256491387e-25
+ uc1 = -7.3692013666e-11 luc1 = 1.67031784950957e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.41 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0191663245768 lvth0 = 2.26029339340689e-8
+ k1 = 0.51047242407276 lk1 = -2.94947323441476e-8
+ k2 = -0.014917698045952 lk2 = 1.70894167977859e-08 wk2 = 6.61744490042422e-24 pk2 = -3.15544362088405e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 69602.3155281761 lvsat = 0.00960414852196073
+ ua = -1.5165106213508e-09 lua = 1.57378335232962e-16
+ ub = 1.5753040065058e-18 lub = -8.05615559377569e-26
+ uc = -5.27318395745652e-11 luc = 2.24839668062795e-17 puc = 4.70197740328915e-38
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00663341319120002 lu0 = 4.34969606879781e-10
+ a0 = 1.113099680712 la0 = -5.32803464830964e-8
+ keta = -0.00348616462015641 lketa = -4.39588448968729e-9
+ a1 = 0.0
+ a2 = 0.75935673367364 la2 = 4.03725008860941e-8
+ ags = 0.277159512155241 lags = 3.57875223277558e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.272911688847361 lvoff = -3.2520436991481e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.2567334619324 lnfactor = 3.19170563265793e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.243261151015 letab = 2.2319990121863e-5
+ dsub = 0.231063940416441 ldsub = 2.87432875546143e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.63111242831704 lpclm = -4.07971696129197e-9
+ pdiblc1 = 0.5605837704226 lpdiblc1 = -1.83253587271965e-7
+ pdiblc2 = 0.000274683463070081 lpdiblc2 = 1.54281818160893e-10
+ pdiblcb = 0.220458260914565 lpdiblcb = -2.1976148752307e-07 wpdiblcb = -2.9778502051909e-23 ppdiblcb = 8.67746995743113e-29
+ drout = 0.522027289967841 ldrout = 2.35802100821845e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.437709665876e-09 lpscbe2 = 1.91688400668287e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.37476536438882 lbeta0 = 4.98971493524157e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.12587401723994e-12 lagidl = 1.05418863444537e-16
+ bgidl = 1394201615.9452 lbgidl = -194.474636807174
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391504383880001 lkt1 = -5.76986497454084e-8
+ kt2 = -0.0452685267320001 lkt2 = -4.89365310308852e-9
+ at = 55827.0751880002 lat = 0.00890619382090246
+ ute = -0.49488123272 lute = 8.74447686476193e-8
+ ua1 = -4.78189710399998e-11 lua1 = 2.97990444514932e-16
+ ub1 = 6.06412088160001e-19 lub1 = -9.32665790686781e-26
+ uc1 = 1.6366545464e-10 luc1 = -6.87444079011884e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.42 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.951579035816 lvth0 = -1.07404439286061e-8
+ k1 = 0.139138830563601 lk1 = 1.53698240010475e-7
+ k2 = 0.117740448063352 lk2 = -4.83558876874859e-08 wk2 = -1.05879118406788e-22 pk2 = -3.78653234506086e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70255.1058400003 lvsat = 0.00928210225510606
+ ua = -4.86169000896802e-10 lua = -3.50928339118575e-16
+ ub = 1.0420180418272e-18 lub = 1.82528675304854e-25
+ uc = -7.86051795167599e-12 luc = 3.47238739486536e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01055413854848 lu0 = -1.49927319943002e-9
+ a0 = 1.49585434488 la0 = -2.42107766994409e-07 wa0 = 3.3881317890172e-21
+ keta = 0.050567389226496 lketa = -3.10625566372871e-08 wketa = -5.29395592033938e-23 pketa = -1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.88128653265272 la2 = -1.97801022826479e-8
+ ags = 1.097940292214 lags = -4.70471251950699e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.26197424659896 lvoff = -3.79162928754222e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.1099157291336 lnfactor = 3.91601329929288e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.681857840994881 leta0 = -9.46507635607321e-8
+ etab = -0.000870723701341264 letab = 1.99713232889716e-10
+ dsub = 0.0824405601279206 ldsub = 1.02064848739392e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.40264312934008 lpclm = 1.08632870057403e-7
+ pdiblc1 = -0.00365505965855961 lpdiblc1 = 9.51068686826147e-8
+ pdiblc2 = -0.00640266916101695 lpdiblc2 = 3.44847360702275e-09 wpdiblc2 = -3.30872245021211e-24 ppdiblc2 = -1.18329135783152e-30
+ pdiblcb = -0.3225732332316 lpdiblcb = 4.81365837360111e-8
+ drout = 1.40305344137712 ldrout = -1.98841578662105e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4174066817368e-09 lpscbe2 = -4.64517597278732e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.8374004106232 lbeta0 = -2.22601954915031e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.08500774325672e-09 lagidl = 1.1310102870514e-15 pagidl = 5.64237288394698e-37
+ bgidl = 1000000000.0
+ cgidl = 532.846726441352 lcgidl = -0.000114872138329124
+ egidl = -1.1321491658048 legidl = 6.07866005159808e-07 wegidl = 8.470329472543e-22 pegidl = -1.0097419586829e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.48341565304 lkt1 = -1.23553280405526e-8
+ kt2 = -0.049672987568 lkt2 = -2.72076520317801e-9
+ at = 91080.1031920002 lat = -0.00848546450853488
+ ute = -0.33479019576 lute = 8.46577665584676e-9
+ ua1 = 9.01049146560001e-10 lua1 = -1.70122254885617e-16 wua1 = 1.57772181044202e-30
+ ub1 = 4.4136286032e-19 lub1 = -1.18415231045482e-26
+ uc1 = 4.74074714316e-11 luc1 = -1.13899269811227e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.43 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.785792300714288 lvth0 = -5.10826564747865e-8
+ k1 = 0.109830032788 lk1 = 1.60830184243594e-7
+ k2 = 0.140327289931343 lk2 = -5.38521246139592e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 199357.877371429 lvsat = -0.0221335079638087
+ ua = -1.20274672320286e-09 lua = -1.76557749328064e-16
+ ub = 1.15786067182572e-18 lub = 1.54339761406273e-25
+ uc = -2.29894954758249e-11 luc = 4.02869387225787e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679047121600002 lu0 = -5.83429918079004e-10
+ a0 = -0.464755997999996 la0 = 2.34983232621324e-7
+ keta = -0.327136074690686 lketa = 6.08470488653921e-8
+ a1 = 0.0
+ a2 = 1.117265914878 la2 = -7.72028531945829e-8
+ ags = 0.04929956616715 lags = 2.0812701179972e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.218487508549716 lvoff = -4.84982687388494e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.36988594933716 lnfactor = 3.28340696485398e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.567449993717428 leta0 = -6.68109868199315e-8
+ etab = 0.193850720008982 letab = -4.71834134366929e-08 wetab = 4.01182597088218e-23 petab = 8.97329279688901e-30
+ dsub = 1.07184049999343 ldsub = -1.38693753827601e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.38934427018857 lpclm = -1.31469012154386e-7
+ pdiblc1 = 0.898253486238859 lpdiblc1 = -1.24361753058971e-7
+ pdiblc2 = 0.0170353361227257 lpdiblc2 = -2.25488372271263e-9
+ pdiblcb = -0.433203011048126 lpdiblcb = 7.50570126103288e-8
+ drout = -0.439476576346854 ldrout = 2.49515990790812e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.60635267050003e-09 lpscbe2 = 1.50908501258468e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.76940471184574 lbeta0 = -2.06056017565909e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.16250109563772e-09 lagidl = -1.36259801878749e-15
+ bgidl = 1000000000.0
+ cgidl = -531.595451576256 lcgidl = 0.000144147092385325
+ egidl = 4.50053273501714 legidl = -7.62779543222403e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.376180031714286 lkt1 = -3.84498296627094e-8
+ kt2 = 0.0904601689714282 lkt2 = -3.68204872491695e-8
+ at = 26226.478514286 lat = 0.00729588681329074
+ ute = -0.3
+ ua1 = 3.68606868285714e-10 lua1 = -4.05588157749091e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -3.26380050227181 lvth0 = 3.78450329166792e-07 wvth0 = 4.32374301974468e-06 pvth0 = -7.49468967556504e-13
+ k1 = -4.6307136029321 lk1 = 9.82546536972046e-07 wk1 = 7.42601738700357e-06 pk1 = -1.28721100182843e-12
+ k2 = 1.02422191607785 lk2 = -2.07064651320942e-07 wk2 = -1.15912305740656e-06 pk2 = 2.00920072524738e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 363519.32933208 lvsat = -0.0505889257237641 wvsat = -0.271997448857645 pvsat = 4.71474937900866e-8
+ ua = 1.03960618389328e-08 lua = -2.18707202787153e-15 wua = -1.93579282067587e-14 pua = 3.35546455950314e-21
+ ub = -3.57142310780033e-18 lub = 9.74104353199095e-25 wub = 6.72394316230623e-24 pub = -1.16551485986784e-30
+ uc = 6.41418596172956e-13 luc = -6.74415111540877e-20 wuc = 6.55503634637616e-19 puc = -1.13623689020815e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.046625333803371 lu0 = -7.48832532924873e-09 wu0 = -6.94985774249307e-08 pu0 = 1.20467444136826e-14
+ a0 = 8.58968829925363 la0 = -1.33449603297603e-06 wa0 = -1.26394969896403e-05 pa0 = 2.19090512919027e-12
+ keta = 2.04794846789243 lketa = -3.5084535557688e-07 wketa = -3.5336991662667e-06 pketa = 6.12524346082338e-13
+ a1 = 0.0
+ a2 = -0.893484834715334 la2 = 2.71336660238426e-7
+ ags = 37.545363627095 lags = -6.29136574039339e-06 wags = -6.27816221301311e-05 pags = 1.08824408167927e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -3.92087664490584 lvoff = 5.93266459378849e-07 wvoff = 5.79962510539864e-06 pvoff = -1.00529541651959e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 41.9938193494667 lnfactor = -6.71333067122626e-06 wnfactor = -7.78511966309952e-05 pnfactor = 1.34945707216235e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.225074950427021 leta0 = -7.46438156605941e-09 weta0 = -1.05802190212116e-06 peta0 = 1.83395400469877e-13
+ etab = -1.36540444630799 letab = 2.23094758582359e-07 wetab = 1.87075980821804e-06 petab = -3.24273763636898e-13
+ dsub = 0.318486163890462 ldsub = -8.10881991618481e-09 wdsub = 1.58254023669715e-08 pdsub = -2.7431435954861e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.354485082557115 lpclm = 1.70802880191845e-07 wpclm = 2.95157094618367e-06 ppclm = -5.11619404669587e-13
+ pdiblc1 = 0.95148729129 lpdiblc1 = -1.33589194358926e-7
+ pdiblc2 = 0.0212117343376134 lpdiblc2 = -2.97881223648482e-9
+ pdiblcb = 0.763376357191859 lpdiblcb = -1.32355661921654e-07 wpdiblcb = -1.3221774355697e-06 ppdiblcb = 2.29183592326781e-13
+ drout = 1.0
+ pscbe1 = 1369148945.55987 lpscbe1 = -98.6551399254558 wpscbe1 = -984.4809492204 ppscbe1 = 0.000170647958775967
+ pscbe2 = 1.09522527291816e-08 lpscbe2 = -2.55725123113284e-16 wpscbe2 = -1.27679985792491e-15 ppscbe2 = 2.21317933772982e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.3849219927818 lbeta0 = -1.35277655200882e-06 wbeta0 = -4.87962787989939e-06 pbeta0 = 8.45824937445994e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.50812115916652e-09 lagidl = -7.29155109359447e-16 wagidl = -7.11547126116867e-15 pagidl = 1.23338155746846e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0640181706666674 lkt1 = -9.25593423329808e-8
+ kt2 = -0.131324749333333 lkt2 = 1.62326691994133e-9
+ at = 615462.065218183 lat = -0.0948410313147893 wat = -0.705986371733274 pat = 1.22374265703502e-7
+ ute = -0.718403621999999 lute = 7.25252470302358e-8
+ ua1 = 8.98188337989136e-10 lua1 = -1.32355408570361e-16 wua1 = -1.56962326948797e-15 pua1 = 2.72075358286506e-22
+ ub1 = 5.46403897747175e-20 lub1 = 5.85985767172297e-26 wub1 = 7.81370639380857e-25 pub1 = -1.35441223888999e-31
+ uc1 = -2.73406652366667e-11 luc1 = 4.84325703289333e-18 wuc1 = 1.23259516440783e-32 puc1 = -2.93873587705572e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.45 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.034517
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29720858
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.911951
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.46 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.034517
+ k1 = 0.42302944
+ k2 = 0.023080264
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -1.9280657e-10
+ ub = 9.7328962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0126711
+ a0 = 1.118778
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17518243
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29720858
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.911951
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.47 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.03968537770652 lvth0 = 4.13125899196556e-8
+ k1 = 0.390669914700908 lk1 = 2.5866062323523e-7
+ k2 = 0.0351772658317135 lk2 = -9.66954244275032e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77014.5327768419 lvsat = -0.188455195353377
+ ua = -9.89907109822339e-11 lua = -7.49901870889346e-16
+ ub = 9.85477846643298e-19 lub = -9.74246151805995e-26
+ uc = -1.11957558265435e-10 luc = 1.06707307552853e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0132665066958 lu0 = -4.75928696699256e-9
+ a0 = 1.126848536098 la0 = -6.45105228724895e-8
+ keta = 0.00968353076963805 lketa = -7.73640015766657e-08 wketa = 7.65142066611551e-24 pketa = -8.36192559534273e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0172899885681765 lags = 1.26208765200977e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.299343388544763 lvoff = 1.70642462635792e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.00110676335524 lnfactor = -7.12652151146605e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.114734399685773 lpclm = 2.1062873248466e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168818489704996 lpdiblc2 = 1.84418379958404e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714327962.849655 lpscbe1 = 342.117401489872
+ pscbe2 = 1.02346458760092e-08 lpscbe2 = -2.88883132878909e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.10658131246379e-11 lalpha0 = -2.59782056161903e-17
+ alpha1 = -8.83803561262885e-13 lalpha1 = 7.06504462287933e-18 walpha1 = 1.85521220424177e-33 palpha1 = -4.32200803793546e-39
+ beta0 = 16.3482835524883 lbeta0 = -5.33042079449266e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.43208327881965e-11 lagidl = 2.85195643082482e-16
+ bgidl = 1704493843.79724 lbgidl = -2813.28203720157
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435787145678042 lkt1 = -6.82083867015442e-8
+ kt2 = -0.0538995747481872 lkt2 = 9.87142670363705e-9
+ at = 133605.523841314 lat = -0.348553690730682
+ ute = -0.186865964192179 lute = 1.24890903956579e-7
+ ua1 = 2.03850284894073e-09 lua1 = 5.70407405815369e-16
+ ub1 = -5.540650054973e-19 lub1 = -1.47404310356667e-24
+ uc1 = 3.51135925346025e-10 luc1 = -1.92270285751065e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0373096643247 lvth0 = 3.18255633950442e-8
+ k1 = 0.397876315328929 lk1 = 2.29883029764097e-7
+ k2 = 0.0322306662092167 lk2 = -8.4928656184203e-08 pk2 = -8.07793566946316e-28
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35013.0233625527 lvsat = -0.0207289717519412
+ ua = 2.2530214708256e-10 lua = -2.04491286412813e-15
+ ub = 7.30246469819167e-19 lub = 9.21800540683505e-25
+ uc = -1.05894772401042e-10 luc = 8.24965543747053e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0145390637694001 lu0 = -9.8410374861681e-9
+ a0 = 1.279695175654 la0 = -6.74878816783818e-7
+ keta = 0.00236686763209581 lketa = -4.8146092636319e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0789146275940666 lags = 1.0159996392514e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.295223607325795 lvoff = 6.12567370160172e-10
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.89071859403239 lnfactor = -2.71834879839183e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.409660780614232 lpclm = 1.22001243377414e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0485835162604493 lpdiblcb = 9.41769516564715e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.98760699558733e-09 lpscbe2 = -1.90232158012228e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.11925577824438e-11 lalpha0 = 1.42773752745155e-16 palpha0 = -1.50463276905253e-36
+ alpha1 = -9.78990408614231e-11 lalpha1 = 3.94479678312631e-16 walpha1 = 2.46519032881566e-31 palpha1 = -2.82118644197349e-37
+ beta0 = -0.505055838463818 lbeta0 = 1.39968726718595e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.12641733093649e-10 lagidl = 9.22339556984973e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431177870254608 lkt1 = -8.66147814024206e-8
+ kt2 = -0.0466701021920688 lkt2 = -1.89983007746662e-8
+ at = 65353.8521233695 lat = -0.0760016964958936
+ ute = 0.732948084020652 lute = -3.54823748770557e-06 wute = -6.7762635780344e-21 pute = 1.29246970711411e-26
+ ua1 = 4.53070332482936e-09 lua1 = -9.38179145816882e-15 wua1 = 5.04870979341448e-29
+ ub1 = -2.45594843985465e-18 lub1 = 6.12082028642299e-24 wub1 = 2.35098870164458e-38
+ uc1 = -2.7031855873761e-10 luc1 = 5.58974949050908e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.49 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.04610950368219 lvth0 = 4.93666175802737e-8
+ k1 = 0.545408083969797 lk1 = -6.41976508749536e-8
+ k2 = -0.0229531449202711 lk2 = 2.50713315250286e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -29678.9552125637 lvsat = 0.108224007437025 pvsat = -8.470329472543e-22
+ ua = -2.46780240508439e-10 lua = -1.1038931018122e-15
+ ub = 8.93180803063207e-19 lub = 5.97017342723471e-25
+ uc = -9.86909462006028e-11 luc = 6.81368938639742e-17 wuc = 1.57772181044202e-30
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0121160398103999 lu0 = -5.01113175378287e-9
+ a0 = 0.823582341107993 la0 = 2.34308228604449e-7
+ keta = -0.0355693011631475 lketa = 2.74735141976551e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.540114866427672 lags = 9.66716775752742e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.284253879441657 lvoff = -2.12538080709266e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.92947467407737 lnfactor = -3.49088846923897e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.327268580000002 leta0 = 8.11823936720047e-7
+ etab = 22.482326763364 letab = -4.49544099258304e-05 wetab = 1.01643953670516e-19 petab = 2.81112161297318e-25
+ dsub = 0.858001399999992 ldsub = -5.94017514673198e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.205964285087447 lpclm = 4.18236089338124e-7
+ pdiblc1 = 0.40380624592791 lpdiblc1 = -2.75205146454694e-8
+ pdiblc2 = 1.43232999999868e-06 lpdiblc2 = 4.2571255218246e-10
+ pdiblcb = -0.00189449793638372 lpdiblcb = 1.10995724841424e-9
+ drout = 0.36191763501607 ldrout = 3.94845105252322e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.06879873224827e-08 lpscbe2 = -3.29841630017526e-15 wpscbe2 = 2.01948391736579e-28
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.19602200021331e-12 lalpha0 = 9.81457458983526e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.17218150587212 lbeta0 = 4.6735577383753e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.17433202659919e-10 lagidl = -1.16650862663801e-16
+ bgidl = 802899192.027405 lbgidl = 392.888530362499
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499503183519998 lkt1 = 4.95806618913848e-8
+ kt2 = -0.0621669880280002 lkt2 = 1.18922306437576e-8
+ at = -10090.7286460004 lat = 0.0743848532457601
+ ute = -1.68308465449999 lute = 1.26773237923172e-6
+ ua1 = -6.01058397519999e-10 lua1 = 8.47544189935723e-16 wua1 = -6.31088724176809e-30 pua1 = 6.01853107621011e-36
+ ub1 = 7.16179343459997e-19 lub1 = -2.02302564913869e-25
+ uc1 = -7.36920136659996e-11 luc1 = 1.67031784950959e-16 wuc1 = -3.94430452610506e-31 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.50 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0191663245768 lvth0 = 2.26029339340765e-8
+ k1 = 0.510472424072759 lk1 = -2.94947323441447e-8
+ k2 = -0.0149176980459521 lk2 = 1.7089416797786e-08 pk2 = -5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 69602.3155281767 lvsat = 0.00960414852196134
+ ua = -1.51651062135081e-09 lua = 1.57378335232956e-16
+ ub = 1.57530400650579e-18 lub = -8.05615559377525e-26
+ uc = -5.27318395745649e-11 luc = 2.24839668062795e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00663341319120003 lu0 = 4.3496960687982e-10
+ a0 = 1.11309968071201 la0 = -5.32803464831032e-8
+ keta = -0.00348616462015638 lketa = -4.39588448968723e-9
+ a1 = 0.0
+ a2 = 0.759356733673641 la2 = 4.03725008861001e-8
+ ags = 0.277159512155237 lags = 3.57875223277557e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.272911688847365 lvoff = -3.25204369914785e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.25673346193241 lnfactor = 3.1917056326579e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.2432611510153 letab = 2.2319990121863e-5
+ dsub = 0.231063940416441 ldsub = 2.87432875546154e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.631112428317024 lpclm = -4.07971696129197e-9
+ pdiblc1 = 0.560583770422603 lpdiblc1 = -1.83253587271961e-7
+ pdiblc2 = 0.00027468346307008 lpdiblc2 = 1.54281818160896e-10
+ pdiblcb = 0.220458260914567 lpdiblcb = -2.1976148752307e-07 wpdiblcb = 5.82335151237331e-22 ppdiblcb = -2.39813715187188e-28
+ drout = 0.522027289967838 ldrout = 2.35802100821851e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.43770966587597e-09 lpscbe2 = 1.91688400668291e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.37476536438874 lbeta0 = 4.98971493524225e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.12587401724014e-12 lagidl = 1.05418863444536e-16
+ bgidl = 1394201615.94521 lbgidl = -194.474636807165
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391504383879997 lkt1 = -5.76986497454101e-8
+ kt2 = -0.0452685267320003 lkt2 = -4.89365310308889e-9
+ at = 55827.0751879988 lat = 0.00890619382090296
+ ute = -0.494881232719997 lute = 8.74447686476193e-8
+ ua1 = -4.78189710399998e-11 lua1 = 2.97990444514927e-16 pua1 = 3.00926553810506e-36
+ ub1 = 6.06412088159995e-19 lub1 = -9.32665790686762e-26
+ uc1 = 1.63665454639999e-10 luc1 = -6.87444079011878e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.951579035815996 lvth0 = -1.07404439286048e-8
+ k1 = 0.13913883056361 lk1 = 1.53698240010471e-7
+ k2 = 0.117740448063352 lk2 = -4.83558876874858e-08 wk2 = 4.2351647362715e-22 pk2 = -2.01948391736579e-28
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70255.1058399994 lvsat = 0.00928210225510595
+ ua = -4.86169000896822e-10 lua = -3.50928339118571e-16
+ ub = 1.04201804182721e-18 lub = 1.82528675304856e-25
+ uc = -7.86051795167597e-12 luc = 3.47238739486555e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0105541385484801 lu0 = -1.49927319943001e-9
+ a0 = 1.49585434488003 la0 = -2.4210776699441e-7
+ keta = 0.0505673892264957 lketa = -3.1062556637287e-08 wketa = -4.2351647362715e-22 pketa = -2.01948391736579e-28
+ a1 = 0.0
+ a2 = 0.881286532652723 la2 = -1.9780102282645e-8
+ ags = 1.09794029221402 lags = -4.70471251950711e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.26197424659896 lvoff = -3.79162928754216e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.10991572913366 lnfactor = 3.91601329929288e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.68185784099488 leta0 = -9.46507635607311e-8
+ etab = -0.000870723701341267 letab = 1.99713232889717e-10
+ dsub = 0.082440560127921 ldsub = 1.02064848739392e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.402643129340092 lpclm = 1.08632870057402e-7
+ pdiblc1 = -0.00365505965856272 lpdiblc1 = 9.51068686826138e-8
+ pdiblc2 = -0.00640266916101692 lpdiblc2 = 3.44847360702274e-09 wpdiblc2 = 5.29395592033938e-23 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.322573233231598 lpdiblcb = 4.81365837360113e-8
+ drout = 1.40305344137712 ldrout = -1.98841578662106e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4174066817369e-09 lpscbe2 = -4.64517597278543e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.83740041062333 lbeta0 = -2.22601954914976e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.0850077432567e-09 lagidl = 1.1310102870514e-15 wagidl = -6.31088724176809e-30 pagidl = 9.02779661431517e-36
+ bgidl = 1000000000.0
+ cgidl = 532.846726441356 lcgidl = -0.000114872138329124
+ egidl = -1.1321491658048 legidl = 6.07866005159807e-07 pegidl = 3.23117426778526e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.483415653040005 lkt1 = -1.23553280405532e-8
+ kt2 = -0.049672987568 lkt2 = -2.72076520317804e-9
+ at = 91080.1031920016 lat = -0.0084854645085346
+ ute = -0.334790195760007 lute = 8.46577665584697e-9
+ ua1 = 9.01049146560002e-10 lua1 = -1.70122254885617e-16 pua1 = -3.00926553810506e-36
+ ub1 = 4.41362860320004e-19 lub1 = -1.18415231045478e-26
+ uc1 = 4.74074714316003e-11 luc1 = -1.13899269811226e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.785792300714292 lvth0 = -5.10826564747874e-8
+ k1 = 0.109830032788011 lk1 = 1.608301842436e-7
+ k2 = 0.140327289931342 lk2 = -5.38521246139583e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 199357.87737143 lvsat = -0.0221335079638085
+ ua = -1.20274672320286e-09 lua = -1.76557749328069e-16
+ ub = 1.15786067182574e-18 lub = 1.54339761406275e-25
+ uc = -2.29894954758248e-11 luc = 4.02869387225789e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679047121599996 lu0 = -5.83429918079021e-10
+ a0 = -0.464755998000015 la0 = 2.34983232621319e-7
+ keta = -0.327136074690687 lketa = 6.08470488653919e-08 wketa = -3.3881317890172e-21
+ a1 = 0.0
+ a2 = 1.11726591487798 la2 = -7.72028531945821e-8
+ ags = 0.04929956616715 lags = 2.08127011799721e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.218487508549714 lvoff = -4.84982687388487e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.36988594933712 lnfactor = 3.28340696485388e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.567449993717432 leta0 = -6.6810986819931e-8
+ etab = 0.193850720008983 letab = -4.71834134366926e-08 wetab = -7.17992771696028e-22 petab = 1.73549399148623e-29
+ dsub = 1.07184049999343 ldsub = -1.386937538276e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.38934427018856 lpclm = -1.31469012154386e-7
+ pdiblc1 = 0.898253486238843 lpdiblc1 = -1.24361753058972e-7
+ pdiblc2 = 0.0170353361227258 lpdiblc2 = -2.25488372271259e-9
+ pdiblcb = -0.433203011048128 lpdiblcb = 7.50570126103286e-8
+ drout = -0.439476576346863 ldrout = 2.49515990790809e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.60635267050024e-09 lpscbe2 = 1.50908501258494e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.76940471184571 lbeta0 = -2.06056017565902e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.16250109563776e-09 lagidl = -1.36259801878749e-15
+ bgidl = 1000000000.0
+ cgidl = -531.595451576264 lcgidl = 0.000144147092385324
+ egidl = 4.50053273501715 legidl = -7.62779543222397e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.376180031714298 lkt1 = -3.84498296627107e-8
+ kt2 = 0.0904601689714273 lkt2 = -3.68204872491697e-8
+ at = 26226.4785142858 lat = 0.00729588681329041
+ ute = -0.3
+ ua1 = 3.68606868285714e-10 lua1 = -4.05588157749085e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.53 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = 4.01114330042014 lvth0 = -8.82573879704224e-07 wvth0 = -8.26003427840006e-06 pvth0 = 1.43177782174931e-12
+ k1 = -0.337578251893376 lk1 = 2.38383041493692e-7
+ k2 = -0.874877798950216 lk2 = 1.22121495082591e-07 wk2 = 2.12582986168546e-06 pk2 = -3.68487096564832e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4323.3989690505 lvsat = 0.0116733784535028 wvsat = 0.34931890995955 pvsat = -6.0550241214568e-8
+ ua = 1.74652235615312e-09 lua = -6.87778153005483e-16 wua = -4.39645475282877e-15 pua = 7.62072673945822e-22
+ ub = 3.02291348007139e-18 lub = -1.68944762269392e-25 wub = -4.68255911473907e-24 pub = 8.11665431830666e-31
+ uc = 1.02037890288087e-12 luc = -1.33129732798224e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0113547034459058 lu0 = -1.37458480434643e-09 wu0 = -8.48947967502222e-09 pu0 = 1.47154942790896e-15
+ a0 = 1.28253178214936 la0 = -6.78881366141971e-8
+ keta = 0.00504336546346629 lketa = 3.26772906795149e-9
+ a1 = 0.0
+ a2 = -0.893484834715338 la2 = 2.71336660238429e-7
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -2.73636761547218 lvoff = 3.87946033234868e-07 wvoff = 3.75072985090612e-06 pvoff = -6.50144010896371e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 49.0978064798815 lnfactor = -7.94472159243803e-06 wnfactor = -9.01392629587307e-05 pnfactor = 1.56245595627403e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.386589552018002 leta0 = 9.85603199587557e-8
+ etab = -0.283879229302801 letab = 3.56253405171125e-8
+ dsub = 0.327635158675349 ldsub = -9.69468837420422e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.35187956888265 lpclm = -1.24974955759423e-7
+ pdiblc1 = 0.951487291290007 lpdiblc1 = -1.33589194358926e-7
+ pdiblc2 = 0.0212117343376135 lpdiblc2 = -2.97881223648482e-9
+ pdiblcb = -0.00100196205692768 lpdiblcb = 1.40147180292528e-10
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.02141081328798e-08 lpscbe2 = -1.27776615079535e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.5639074624669 lbeta0 = -8.63787535353047e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.94518992804005e-10 lagidl = -1.61115370464976e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0640181706666567 lkt1 = -9.25593423329778e-8
+ kt2 = -0.131324749333331 lkt2 = 1.62326691994176e-9
+ at = 207316.636533339 lat = -0.0240939189974152
+ ute = -0.718403622000011 lute = 7.25252470302352e-8
+ ua1 = -9.24357266666552e-12 lua1 = 2.4937023958895e-17
+ ub1 = 5.0636703399999e-19 lub1 = -1.97028163394924e-26
+ uc1 = -2.73406652366669e-11 luc1 = 4.84325703289333e-18 puc1 = 1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.54 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.13241955778733 wvth0 = 1.66409108959069e-7
+ k1 = 0.192177033644933 wk1 = 3.92389577053255e-7
+ k2 = 0.10889696070478 wk2 = -1.45866260853715e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47393.65057134 wvsat = 0.0102738357954393
+ ua = 3.84222479981006e-09 wua = -6.85851309758997e-15
+ ub = -1.01712351918573e-18 wub = 3.38318920810846e-24
+ uc = -2.9907055997136e-10 wuc = 3.40734625110569e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0309163958791707 wu0 = -3.10122993573125e-8
+ a0 = 0.68344991754 wa0 = 7.3994551260234e-7
+ keta = -0.0222783333676765 wketa = 3.78758723671381e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.0822918634785329 wags = 4.37639922040647e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.289281852289933 wvoff = -1.347339359671e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.381769632056 wnfactor = -7.98570555251856e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.642546162609021 wpclm = -8.39290566185525e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00107066232286653 wpdiblc2 = 2.14601346288427e-9
+ pdiblcb = 0.646662666666666 wpdiblcb = -1.14165337869787e-6
+ drout = 0.56
+ pscbe1 = 613201011.8902 wpscbe1 = 244.639251336941
+ pscbe2 = 6.85502405793333e-09 wpscbe2 = 5.13019070518567e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.76469737917133e-11 walpha0 = -1.01697518277301e-16
+ alpha1 = 2.7482008494454e-16 walpha1 = -3.59943462659449e-22
+ beta0 = -58.562215686586 wbeta0 = 0.000115993671210224
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.68598976745332e-11 wagidl = 2.66621387565086e-16
+ bgidl = 2536481961.69 wbgidl = -2012.39526476418
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.104157749960667 wkt1 = -5.78188641161467e-7
+ kt2 = -0.05327118983764 wkt2 = 1.03101574976824e-9
+ at = 358665.066666667 wat = -0.456661351479146
+ ute = 3.48347113841513 wute = -6.21206945336434e-6
+ ua1 = 1.00553410450693e-08 wua1 = -1.35052639924294e-14
+ ub1 = -4.87864951938746e-18 wub1 = 7.03723111369948e-24
+ uc1 = 4.544979784468e-10 wuc1 = -5.84541713883244e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.55 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.13241955778733 wvth0 = 1.66409108959069e-7
+ k1 = 0.192177033644934 wk1 = 3.92389577053254e-7
+ k2 = 0.10889696070478 wk2 = -1.45866260853715e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47393.65057134 wvsat = 0.0102738357954394
+ ua = 3.84222479981006e-09 wua = -6.85851309758997e-15
+ ub = -1.01712351918573e-18 wub = 3.38318920810846e-24
+ uc = -2.9907055997136e-10 wuc = 3.4073462511057e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0309163958791707 wu0 = -3.10122993573125e-8
+ a0 = 0.683449917539999 wa0 = 7.39945512602341e-7
+ keta = -0.0222783333676765 wketa = 3.78758723671381e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.0822918634785332 wags = 4.37639922040648e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.289281852289933 wvoff = -1.347339359671e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.381769632056 wnfactor = -7.98570555251856e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.642546162609021 wpclm = -8.39290566185525e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00107066232286653 wpdiblc2 = 2.14601346288427e-9
+ pdiblcb = 0.646662666666666 wpdiblcb = -1.14165337869787e-6
+ drout = 0.56
+ pscbe1 = 613201011.8902 wpscbe1 = 244.639251336941
+ pscbe2 = 6.85502405793333e-09 wpscbe2 = 5.13019070518566e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.76469737917133e-11 walpha0 = -1.01697518277301e-16
+ alpha1 = 2.7482008494454e-16 walpha1 = -3.59943462659448e-22
+ beta0 = -58.562215686586 wbeta0 = 0.000115993671210224
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.68598976745332e-11 wagidl = 2.66621387565086e-16
+ bgidl = 2536481961.69 wbgidl = -2012.39526476418
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.104157749960666 wkt1 = -5.78188641161466e-7
+ kt2 = -0.05327118983764 wkt2 = 1.03101574976829e-9
+ at = 358665.066666667 wat = -0.456661351479146
+ ute = 3.48347113841513 wute = -6.21206945336434e-6
+ ua1 = 1.00553410450693e-08 wua1 = -1.35052639924294e-14
+ ub1 = -4.87864951938746e-18 wub1 = 7.03723111369948e-24
+ uc1 = 4.544979784468e-10 wuc1 = -5.84541713883244e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.56 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.14806250351302 lvth0 = 1.25039352501092e-07 wvth0 = 1.84213174248057e-07 pvth0 = -1.42313911628938e-13
+ k1 = -0.089708682303987 lk1 = 2.25320780495171e-06 wk1 = 8.16519773306009e-07 pk1 = -3.3902160146546e-12
+ k2 = 0.204376147370209 lk2 = -7.63197410981866e-07 wk2 = -2.87594479143781e-07 pk2 = 1.13288155293028e-12
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 108265.231128122 lvsat = -0.486567117984583 wvsat = -0.0531181307671393 pvsat = 5.06713415219389e-7
+ ua = 6.15438713277867e-09 lua = -1.84818950382866e-14 wua = -1.06291302135854e-14 pua = 3.01398170767368e-20
+ ub = -1.92887118191961e-18 lub = 7.28790723894186e-24 wub = 4.95364202937741e-24 pub = -1.25531602134563e-29
+ uc = -4.09735559396951e-10 luc = 8.84582745178557e-16 wuc = 5.06145834754887e-16 puc = -1.32218770767589e-21
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0421160363720325 lu0 = -8.95225119379315e-08 wu0 = -4.90367630408447e-08 pu0 = 1.44075630491199e-13
+ a0 = 0.471748982998644 la0 = 1.69219712470496e-06 wa0 = 1.11350035560412e-06 pa0 = -2.98595012165015e-12
+ keta = 0.00844478630403462 lketa = -2.45580279950436e-07 wketa = 2.10554624320277e-09 pketa = 2.85924307078845e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.595762931923631 lags = 4.1043478033028e-06 wags = 1.04203191979317e-06 pags = -4.83110952253113e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.235768414400914 lvoff = -4.27750996588934e-07 wvoff = -1.08061066416212e-07 pvoff = 7.56071239479694e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 3.81134522329346 lnfactor = -1.14270808973109e-05 wnfactor = -3.07693870241999e-06 pnfactor = 1.82117666887487e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.384311688958626 lpclm = 8.20802188553403e-06 wpclm = 4.58211894738672e-07 ppclm = -1.03713757259989e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00040472403201286 lpdiblc2 = -1.17932618151389e-08 wpdiblc2 = -4.00978605474555e-10 ppdiblc2 = 2.03589684857112e-14
+ pdiblcb = 0.646662666666666 wpdiblcb = -1.14165337869787e-6
+ drout = 0.56
+ pscbe1 = 426713070.440696 lpscbe1 = 1490.6611489301 wpscbe1 = 488.871169975975 ppscbe1 = -0.0019522282760703
+ pscbe2 = 4.17523356151092e-09 lpscbe2 = 2.14204712070922e-14 wpscbe2 = 1.02994388181522e-14 ppscbe2 = -4.13195473728039e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.18114142186181e-11 lalpha0 = -1.13221159913114e-16 walpha0 = -1.20249283643804e-16 palpha0 = 1.48290531071154e-22
+ alpha1 = -3.85189284509951e-12 lalpha1 = 3.07916781804902e-17 walpha1 = 5.04498660910489e-18 palpha1 = -4.03291603218072e-23
+ beta0 = -29.498457816076 lbeta0 = -0.000232316440209147 wbeta0 = 7.79276410366345e-05 pbeta0 = 3.04274645495696e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.76249913515058e-10 lagidl = 9.54324750438669e-16 wagidl = 4.08908249577133e-16 pagidl = -1.13734698102165e-21
+ bgidl = 4070404912.6728 lbgidl = -12261.164613163 wbgidl = -4021.43888521489 pbgidl = 0.0160589647150062
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.215767293164757 lkt1 = -2.55726900436609e-06 wkt1 = -1.10747457529843e-06 pkt1 = 4.2307613702025e-12
+ kt2 = 0.0276522015489231 lkt2 = -6.46848019459088e-07 wkt2 = -1.38616995657157e-07 pkt2 = 1.11625375620341e-12
+ at = 700484.210779479 lat = -2.73227595376442 wat = -0.963547626469386 pat = 4.05171332355793e-6
+ ute = 7.40343573436436 lute = -3.13336019634556e-05 wute = -1.29015561077682e-05 pute = 5.34713278751395e-11
+ ua1 = 1.70386756795036e-08 lua1 = -5.58201541001395e-14 wua1 = -2.54964267674012e-14 pua1 = 9.58494170733675e-20
+ ub1 = -9.13700837332206e-18 lub1 = 3.40385016447918e-23 wub1 = 1.45887910425019e-23 pub1 = -6.03621709381733e-29
+ uc1 = 1.20714519046778e-09 luc1 = -6.01616356044138e-15 wuc1 = -1.45499507151844e-15 puc1 = 6.95782790081299e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.57 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.13309937680618 lvth0 = 6.52865300238187e-08 wvth0 = 1.6281781663063e-07 pvth0 = -5.68750170316811e-14
+ k1 = 0.262056531028444 lk1 = 8.4849041147321e-07 wk1 = 2.30858618970434e-07 pk1 = -1.05147307192248e-12
+ k2 = 0.0957324515871884 lk2 = -3.29346412151091e-07 wk2 = -1.07936664382282e-07 pk2 = 4.15447174246221e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 44830.6131584935 lvsat = -0.233251247530985 wvsat = -0.0166873716784494 pvsat = 3.61233080581679e-7
+ ua = 3.09892228816686e-09 lua = -6.28039116663418e-15 wua = -4.88441342057092e-15 pua = 7.19922120795389e-21
+ ub = -6.0803066611114e-19 lub = 2.01334461522432e-24 wub = 2.27472612323588e-24 pub = -1.85534352665691e-30
+ uc = -2.4633154526909e-10 luc = 2.32055286209232e-16 wuc = 2.38706309275638e-16 puc = -2.54211287877633e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0281504448662749 lu0 = -3.37531846855121e-08 wu0 = -2.31358388506404e-08 pu0 = 4.06444856873366e-14
+ a0 = 1.4963528413622 la0 = -2.39939239784484e-06 wa0 = -3.68262177357714e-07 pa0 = 2.9312285082026e-12
+ keta = -0.0274058270029605 lketa = -1.02416663508307e-07 wketa = 5.06059054789188e-08 pketa = 9.22459795292096e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.434971147811929 lags = 3.46225186172174e-06 wags = 8.73473338437298e-07 pags = -4.15799813437665e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.345784949781473 lvoff = 1.15822147745914e-08 wvoff = 8.59412474605751e-08 pvoff = -1.86455726124082e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.211017464811619 lnfactor = 2.95024475308949e-06 wnfactor = 2.85505889272422e-06 pnfactor = -5.47670472384933e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.18609657993379 leta0 = 1.06261358431964e-06 weta0 = 4.52295586189136e-07 peta0 = -1.80616915156135e-12
+ etab = 0.162625307030371 letab = -9.28951478326047e-07 wetab = -3.95403051147478e-07 petab = 1.57897802946317e-12
+ dsub = -0.444138037485999 ldsub = 4.00986258233826e-06 wdsub = 1.70677579694013e-06 pdsub = -6.81573264740132e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.70974964528105 lpclm = -4.14761081481598e-06 wpclm = -3.90955810702429e-06 ppclm = 7.0706061973012e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00530281481429438 lpdiblc2 = 1.09988699462959e-08 wpdiblc2 = 9.37886269164132e-09 ppdiblc2 = -1.86952434000309e-14
+ pdiblcb = 0.543878313301866 lpdiblcb = 4.10452664097085e-07 wpdiblcb = -1.00703237359627e-06 ppdiblcb = -5.37587175270378e-13
+ drout = 0.56
+ pscbe1 = 800000134.108803 lpscbe1 = -0.000267324172455119 wpscbe1 = -0.000227950391490594 ppscbe1 = 4.54382177716983e-10
+ pscbe2 = 1.11778463431706e-08 lpscbe2 = -6.54332851319534e-15 wpscbe2 = -2.02310004718823e-15 ppscbe2 = 7.888515334637e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.21584610756616e-11 lalpha0 = 5.81499353954794e-16 walpha0 = 1.03626318588601e-16 palpha0 = -7.45720418596394e-22
+ alpha1 = -4.26684481638701e-10 lalpha1 = 1.71930512264835e-15 walpha1 = 5.58850488434739e-16 palpha1 = -2.25186171537118e-21
+ beta0 = -193.323014968594 lbeta0 = 0.000421890389201177 wbeta0 = 0.000327740822051358 pbeta0 = -6.93313823151279e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.66332297459237e-10 lagidl = -8.13055610769002e-16 wagidl = -2.61234337994005e-16 pagidl = 1.5387588793445e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.362519145179734 lkt1 = -2.47975795240377e-07 wkt1 = -1.16702132407964e-07 pkt1 = 2.74272124655165e-13
+ kt2 = -0.176477384525888 lkt2 = 1.68310413537728e-07 wkt2 = 2.20638915650107e-07 pkt2 = -3.1837652614452e-13
+ at = -60799.1601499153 lat = 0.307785860136025 wat = 0.214427598618021 pat = -6.52339905842163e-7
+ ute = 0.667952381135571 lute = -4.43654034063966e-06 wute = 1.1047593901243e-07 pute = 1.50988584551249e-12
+ ua1 = 6.36131383769795e-09 lua1 = -1.31818393175071e-14 wua1 = -3.11156594048633e-15 pua1 = 6.45910170853693e-21
+ ub1 = -1.39515228047283e-18 lub1 = 3.12265351868547e-24 wub1 = -1.80307999769919e-24 pub1 = 5.09611057776103e-30
+ uc1 = -4.34624422706946e-10 luc1 = 5.39977423094566e-16 wuc1 = 2.79277610696139e-16 puc1 = 3.22908965635936e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.58 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.17820063689786 lvth0 = 1.55188585612456e-07 wvth0 = 2.24520873372474e-07 pvth0 = -1.79870064751356e-13
+ k1 = 0.802645567049158 lk1 = -2.29086256410248e-07 wk1 = -4.37237405411771e-07 pk1 = 2.80268121127493e-13
+ k2 = -0.11509478885164 lk2 = 9.09035376507616e-08 wk2 = 1.5661704056752e-07 pk2 = -1.11897778871007e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -390963.785139197 lvsat = 0.635434286782936 wvsat = 0.614091071646121 pvsat = -8.96121560078033e-7
+ ua = 3.29318691110069e-09 lua = -6.66762622158385e-15 wua = -6.01703155420386e-15 pua = 9.45691197321352e-21
+ ub = -1.65175280460187e-18 lub = 4.09383561531915e-24 wub = 4.32573104914663e-24 pub = -5.94368958366198e-30
+ uc = -2.91060830445357e-10 luc = 3.21215870063922e-16 wuc = 3.26979210259922e-16 puc = -4.30169015779845e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0236734912505302 lu0 = -2.48291029190109e-08 wu0 = -1.964468793724e-08 pu0 = 3.36854419079208e-14
+ a0 = -1.88878507956812 la0 = 4.34833165518654e-06 wa0 = 4.61032536682835e-06 pa0 = -6.99277922995015e-12
+ keta = -0.249028955554392 lketa = 3.39353140312146e-07 wketa = 3.62826382566213e-07 pketa = -5.30114961827023e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 3.67528159780154 lags = -4.7308711257139e-06 wags = -5.32897519735221e-06 pags = 8.20557822505693e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.269419496643836 lvoff = -1.40639944851877e-07 wvoff = -2.52146264524148e-08 pvoff = 2.02925654781564e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 3.38072621933057 lnfactor = -3.36805615622581e-06 wnfactor = -2.46675349428202e-06 pnfactor = 5.13146613604091e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.16281092259415 leta0 = 3.00953539868956e-06 weta0 = 1.42020657959414e-06 peta0 = -3.7355429153333e-12
+ etab = 97.9650200521429 letab = -0.000195882181414759 wetab = -0.000128301119152594 petab = 2.56538302351689e-10
+ dsub = 3.867059549944 ldsub = -4.58381139419427e-06 wdsub = -5.11462311971374e-06 pdsub = 6.78162102632368e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.221754719860793 lpclm = 1.69586823338714e-06 wpclm = 7.27012042452521e-07 ppclm = -2.1716452713166e-12
+ pdiblc1 = 0.42428281429169 lpdiblc1 = -6.83372364745678e-08 wpdiblc1 = -3.48048873590841e-08 ppdiblc1 = 6.93779045585817e-14
+ pdiblc2 = -0.000715794823729934 lpdiblc2 = 1.85538869234418e-09 wpdiblc2 = 1.21910126018066e-09 ppdiblc2 = -2.43008086776599e-15
+ pdiblcb = 1.41455173436522 lpdiblcb = -1.3250937516985e-06 wpdiblcb = -2.40759343507404e-06 ppdiblcb = 2.25420440989358e-12
+ drout = 0.868453341004798 ldrout = -6.14851765851821e-07 wdrout = -8.60980115275817e-07 pdrout = 1.71622438102367e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 1.18969441836019e-08 lpscbe2 = -7.97673356424496e-15 wpscbe2 = -2.05491499482408e-15 ppscbe2 = 7.95193327872753e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.18395971471157e-10 lalpha0 = -2.16941017509216e-16 walpha0 = -5.3915813995363e-16 palpha0 = 5.35566268425259e-22
+ alpha1 = 7.69444931387629e-10 lalpha1 = -6.64985089254725e-16 walpha1 = -1.13788380045566e-15 palpha1 = 1.13030321857702e-21
+ beta0 = 27.7942051024633 lbeta0 = -1.88709680208248e-05 wbeta0 = -4.01513503565217e-05 pbeta0 = 4.00196240118995e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.81499121616201e-10 lagidl = 4.78291374467994e-16 wagidl = 1.01803054651621e-15 pagidl = -1.01124842701532e-21
+ bgidl = 140972920.602244 lbgidl = 1712.33132039256 wbgidl = 1125.10401682999 pbgidl = -0.00224271259069986
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.738360763569044 lkt1 = 5.01203584676532e-07 wkt1 = 4.05996308599238e-07 pkt1 = -7.67642540345248e-13
+ kt2 = -0.179245092622563 lkt2 = 1.73827391259737e-07 wkt2 = 1.99002595075393e-07 pkt2 = -2.75248026162759e-13
+ at = -17354.309577376 lat = 0.221185588585461 wat = 0.0123462150321751 pat = -2.4952340484792e-7
+ ute = -5.3249347975136 lute = 7.50930940227453e-06 wute = 6.19020637415626e-06 pute = -1.06090718606162e-11
+ ua1 = -2.39547311000422e-09 lua1 = 4.2733968632517e-15 wua1 = 3.0500424111103e-15 pua1 = -5.82306635981799e-21
+ ub1 = -2.76214515581494e-19 lub1 = 8.92232352292501e-25 wub1 = 1.68681372123368e-24 pub1 = -1.86042718814917e-30
+ uc1 = -5.77073994705279e-10 luc1 = 8.2392756804258e-16 wuc1 = 8.55619595892063e-16 puc1 = -1.11655348352288e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.59 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.01004200544915 lvth0 = -1.18497730335388e-08 wvth0 = -1.55089902675302e-08 pvth0 = 5.85607199370768e-14
+ k1 = 0.885348114424805 lk1 = -3.11237839415278e-07 wk1 = -6.37192030645503e-07 pk1 = 4.78890648647919e-13
+ k2 = -0.146932329533757 lk2 = 1.22528976636855e-07 wk2 = 2.24390840157271e-07 pk2 = -1.79220069407891e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 346418.317349862 lvsat = -0.0970353761393405 wvsat = -0.470515839931597 pvsat = 1.81259700254754e-7
+ ua = -5.38320252327834e-09 lua = 1.95096110638335e-15 wua = 6.5723794001045e-15 pua = -3.04862832531725e-21
+ ub = 3.54116292643623e-18 lub = -1.06448491111878e-24 wub = -3.34145336545218e-24 pub = 1.67241604836677e-30
+ uc = 2.27378112630769e-11 luc = 9.50775490654963e-18 wuc = -1.28278950348005e-16 puc = 2.2056214962113e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0105184400572399 lu0 = 9.13504174238687e-09 wu0 = 2.91537287745804e-08 pu0 = -1.47878797517655e-14
+ a0 = 4.3839777211127 la0 = -1.88264199971615e-06 wa0 = -5.55964943632238e-06 pa0 = 3.10944320106198e-12
+ keta = 0.126745361892265 lketa = -3.39177686316813e-08 wketa = -2.21360021383582e-07 pketa = 5.0179592299658e-14
+ a1 = 0.0
+ a2 = 0.622863910459608 la2 = 1.75956008911874e-07 wa2 = 2.32002611614032e-07 pa2 = -2.30457010215458e-13
+ ags = -2.12186353869076 lags = 1.02765342987908e-06 wags = 4.07772071829569e-06 pags = -1.13845028240093e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.359410493563707 lvoff = -5.12484679534861e-08 wvoff = 1.47025668625934e-07 pvoff = 3.18328245490271e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -0.988608471007618 lnfactor = 9.72170026405347e-07 wnfactor = 3.81650243684772e-06 pnfactor = -1.10993074407564e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 3.22547100492347 leta0 = -1.34951179462693e-06 weta0 = -4.64959550394482e-06 peta0 = 2.29382214672513e-12
+ etab = -197.137625864247 letab = 9.72544906745357e-05 wetab = 0.000258181261645271 petab = -1.27369332825301e-10
+ dsub = -1.67741657416397 ldsub = 9.23727429974888e-07 wdsub = 3.24392486851004e-06 pdsub = -1.52124231520255e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.347851242867 lpclm = -8.5661901441696e-07 wpclm = -2.91801340946853e-06 ppclm = 1.44909702104375e-12
+ pdiblc1 = 0.407050002259573 lpdiblc1 = -5.12192294362095e-08 wpdiblc1 = 2.60967824871713e-07 ppdiblc1 = -2.24424369863334e-13
+ pdiblc2 = 0.00152615705793975 lpdiblc2 = -3.71627305889825e-10 wpdiblc2 = -2.12718248138569e-09 ppdiblc2 = 8.93909931514041e-16
+ pdiblcb = 1.04478401132076 lpdiblcb = -9.57789421224963e-07 wpdiblcb = -1.40114126451208e-06 ppdiblcb = 1.25445722369191e-12
+ drout = -0.491044122009595 ldrout = 7.3558872506397e-07 wdrout = 1.72196023055163e-06 pdrout = -8.49508416219882e-13
+ pscbe1 = 800000000.0
+ pscbe2 = -1.5373240883963e-09 lpscbe2 = 5.36803561252522e-15 wpscbe2 = 1.1855759218561e-14 ppscbe2 = -5.86606802304801e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.04102368697252 lbeta0 = 1.743955700076e-06 wbeta0 = 2.26701701300324e-06 pbeta0 = -2.11615219420968e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.59851478234573e-10 lagidl = -4.56787947686574e-16 wagidl = -9.62015589866671e-16 pagidl = 9.5560664200698e-22
+ bgidl = 2718054158.79551 lbgidl = -847.58140259186 wbgidl = -2250.20803365998 pbgidl = 0.00111011313090975
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.0372088399887707 lkt1 = -2.69199174182381e-07 wkt1 = -7.28701958307797e-07 pkt1 = 3.59496366707652e-13
+ kt2 = 0.0460055339764513 lkt2 = -4.99226156648746e-08 wkt2 = -1.55142372751517e-07 pkt2 = 7.65376278884877e-14
+ at = 305573.687518636 lat = -0.0995910621938978 wat = -0.424504856285423 pat = 1.8441736463256e-7
+ ute = 5.00824121046288 lute = -2.75502698713682e-06 wute = -9.35388944844504e-06 pute = 4.8314691956149e-12
+ ua1 = 3.23896573225266e-09 lua1 = -1.32350534743806e-15 wua1 = -5.58668666250101e-15 pua1 = 2.75612482470492e-21
+ ub1 = 1.26843189565092e-18 lub1 = -6.42123624548278e-25 wub1 = -1.12526300402819e-24 pub1 = 9.32915481968996e-31
+ uc1 = 4.77400120260054e-10 luc1 = -2.23521640368855e-16 wuc1 = -5.33268050757295e-16 puc1 = 2.63081393624503e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.60 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.960607295430903 lvth0 = -3.62377940045217e-08 wvth0 = 1.53457138600076e-08 pvth0 = 4.33389219122074e-14
+ k1 = -0.870839999532857 lk1 = 5.55156492348367e-07 wk1 = 1.71670363862158e-06 pk1 = -6.82375533036964e-13
+ k2 = 0.496158449118115 lk2 = -1.94732141921703e-07 wk2 = -6.43213045632426e-07 pk2 = 2.48801896399827e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 202824.348665743 lvsat = -0.0261950148166546 wvsat = -0.225333536452963 pvsat = 6.03019530212122e-8
+ ua = 2.99483138063512e-10 lua = -8.52523672411721e-16 wua = -1.33540609511111e-15 pua = 8.52582755321427e-22
+ ub = 6.31707987743998e-19 lub = 3.7085976942577e-25 wub = 6.97421314009498e-25 pub = -3.20114308249495e-31
+ uc = 1.1037409937167e-10 luc = -3.37265561963678e-17 wuc = -2.00968368565343e-16 puc = 5.79166671666178e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.015263691195774 lu0 = -3.58426332571251e-09 wu0 = -8.00502537772731e-09 pu0 = 3.54394570422566e-15
+ a0 = 1.65025854981243 la0 = -5.33994451185211e-07 wa0 = -2.62447342981096e-07 pa0 = 4.96132114737178e-13
+ keta = 0.408858957758571 lketa = -1.73095125789173e-07 wketa = -6.0900329893816e-07 pketa = 2.41418751561879e-13
+ a1 = 0.0
+ a2 = 0.251172969660389 la2 = 3.5932527426388e-07 wa2 = 1.07103061381042e-06 pa2 = -6.44381406763023e-13
+ ags = -2.53523781434261 lags = 1.23158666828061e-06 wags = 6.17546614783037e-06 pags = -2.17334781711671e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.521949906309723 lvoff = 2.89384008518076e-08 wvoff = 4.41891599783223e-07 pvoff = -1.13635744196248e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.282152463094171 lnfactor = 3.45255368697438e-07 wnfactor = 1.40698415489704e-06 pnfactor = 7.877618610534e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.32617658651253 leta0 = -4.1251768483692e-07 weta0 = -1.09517576200741e-06 peta0 = 5.40291820077214e-13
+ etab = -0.00395776844010065 letab = 9.61123486551509e-10 wetab = 5.2471802157573e-09 petab = -1.29420113966165e-15
+ dsub = 0.308547421412642 ldsub = -5.60240756748854e-08 wdsub = -3.84323373835187e-07 pdsub = 2.68710416179558e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.31250524601823 lpclm = 4.558359350967e-07 wpclm = 1.21556787285796e-06 ppclm = -5.90155701616637e-13
+ pdiblc1 = 0.465892152337624 lpdiblc1 = -8.02482980714149e-08 wpdiblc1 = -7.9810921112226e-07 ppdiblc1 = 2.98058576919861e-13
+ pdiblc2 = 0.00474571276608955 lpdiblc2 = -1.95995647983704e-09 wpdiblc2 = -1.89493752232203e-08 ppdiblc2 = 9.19293685438523e-15
+ pdiblcb = -1.97568158996172 lpdiblcb = 5.32321037580538e-07 wpdiblcb = 2.80985803510685e-06 ppdiblcb = -8.22988748783494e-13
+ drout = 0.898895496875351 ldrout = 4.98786933625088e-08 wdrout = 8.56938533734916e-07 pdrout = -4.22760342355716e-13
+ pscbe1 = 799767456.074087 lpscbe1 = 0.114722755322418 wpscbe1 = 0.395264724227673 ppscbe1 = -1.94999108521412e-7
+ pscbe2 = 9.40276673535493e-09 lpscbe2 = -2.91269142825731e-17 wpscbe2 = 2.48841346709769e-17 ppscbe2 = -2.94477709118472e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.396648879577 lbeta0 = -1.39151572119309e-06 wbeta0 = -6.04980482296609e-06 pbeta0 = 1.98685205670376e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.12677109608235e-08 lagidl = 5.37819805087344e-15 wagidl = 1.5608228168974e-14 pagidl = -7.21912427349195e-21
+ bgidl = 1906629732.22925 lbgidl = -447.274898838516 wbgidl = -1541.03681564476 pbgidl = 0.000760252020556555
+ cgidl = 1314.81899247236 lcgidl = -0.000500648772108331 wcgidl = -0.00132915125980254 pcgidl = 6.55720824208464e-10
+ egidl = -5.2700921379826 legidl = 2.64927051516806e-06 wegidl = 7.03343629100403e-06 pegidl = -3.46986139293135e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.411109332528258 lkt1 = -4.80267835891742e-08 wkt1 = -1.22902104300533e-07 pkt1 = 6.06322783314164e-14
+ kt2 = 0.0917427465178488 lkt2 = -7.24865206256225e-08 wkt2 = -2.40370290969696e-07 pkt2 = 1.18583798606408e-13
+ at = 183751.546951822 lat = -0.0394915710109467 wat = -0.157517563693496 pat = 5.27023876798438e-8
+ ute = -0.470047706110753 lute = -5.23788896122136e-08 wute = 2.29902898210111e-07 pute = 1.03420246900739e-13
+ ua1 = 1.5568073272951e-09 lua1 = -4.93632684253113e-16 wua1 = -1.11461985279068e-15 pua1 = 5.49884328936051e-22
+ ub1 = -2.96320798163869e-19 lub1 = 1.29828339912921e-25 wub1 = 1.25387204457542e-24 pub1 = -2.40802244639012e-31
+ uc1 = 4.73155848733005e-11 luc1 = -1.13445958502243e-17 wuc1 = 1.5618346075442e-19 puc1 = -7.70512361616663e-26
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.61 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.878886907244986 lvth0 = -5.61234698249064e-08 wvth0 = 1.58236831312625e-07 pvth0 = 8.5680831735206e-15
+ k1 = 3.09060327611239 lk1 = -4.08813191460595e-07 wk1 = -5.06654607030933e-06 pk1 = 9.68246884634865e-13
+ k2 = -0.941669914875341 lk2 = 1.55146136515737e-07 wk2 = 1.83911630929196e-06 pk2 = -3.55243164168764e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 70301.0671297982 lvsat = 0.00605293546573915 wvsat = 0.219363306565091 pvsat = -4.79096873651152e-8
+ ua = -5.60992647605409e-09 lua = 5.85460244268429e-16 wua = 7.49106940890682e-15 pua = -1.29523414087529e-21
+ ub = 3.80296353054249e-18 lub = -4.00827211847729e-25 wub = -4.49599295230153e-24 pub = 9.436407324861e-31
+ uc = -9.89370266206271e-11 luc = 1.7206794580346e-17 wuc = 1.29091223672635e-16 puc = -2.23993738893872e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00607121728030889 lu0 = 1.60733063304055e-09 wu0 = 2.18615547004308e-08 pu0 = -3.72372815883316e-15
+ a0 = -2.46687383977989 la0 = 4.67860310233404e-07 wa0 = 3.4030841850462e-06 pa0 = -3.95830996229929e-13
+ keta = -1.08381757113888 lketa = 1.90129795399675e-07 wketa = 1.28616347147215e-06 pketa = -2.19747340016225e-13
+ a1 = 0.0
+ a2 = 4.4666105048153 la2 = -6.66450864665647e-07 wa2 = -5.69302234185812e-06 pa2 = 1.00156971136345e-12
+ ags = 5.68563527163015 lags = -7.68864146713827e-07 wags = -9.58031765194225e-06 pags = 1.66063310115236e-12
+ b0 = 0.0
+ b1 = 1.75247592434801e-23 lb1 = -4.26443986478995e-30 wb1 = -2.97875728309831e-29 pb1 = 7.24844839754578e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.212808651804103 lvoff = -4.62874137370809e-08 wvoff = -9.6525924582703e-09 pvoff = -3.75788354458727e-15
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 3.03855510498472 lnfactor = -3.25482137374923e-07 wnfactor = -2.83630738169255e-06 pnfactor = 1.11133026203598e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.48955334860311 leta0 = 2.72656406114251e-07 weta0 = 3.49637538648327e-06 peta0 = -5.77007053294212e-13
+ etab = 0.583180912759274 letab = -1.41912028919142e-07 wetab = -6.61760958351805e-07 petab = 1.61014225283092e-13
+ dsub = -0.419015932804587 ldsub = 1.21019735813627e-07 wdsub = 2.53407159296825e-06 pdsub = -4.41445978252457e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.78991247095034 lpclm = -5.42438187314997e-07 wpclm = -4.08034707481284e-06 ppclm = 6.98541649919682e-13
+ pdiblc1 = -0.212048977222925 lpdiblc1 = 8.47205405135901e-08 wpdiblc1 = 1.88722795190995e-06 ppdiblc1 = -3.55385997658071e-13
+ pdiblc2 = -0.0357092232155182 lpdiblc2 = 7.88426673205544e-09 wpdiblc2 = 8.96521533276172e-08 ppdiblc2 = -1.72339419001185e-14
+ pdiblcb = 0.114993147851663 lpdiblcb = 2.35804282305033e-08 wpdiblcb = -9.31792145159875e-07 ppdiblcb = 8.74969227822502e-14
+ drout = 1.36108751115946 ldrout = -6.25901870093584e-08 wdrout = -3.06049476333898e-06 pdrout = 5.30500041287652e-13
+ pscbe1 = 800830514.021122 lpscbe1 = -0.143959639392961 wpscbe1 = -1.4116597293887 ppscbe1 = 2.44694274172813e-7
+ pscbe2 = 8.06601424215027e-09 lpscbe2 = 2.96155763908869e-16 wpscbe2 = 9.18436028947751e-16 ppscbe2 = -2.46882901761371e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.20416726554275 lbeta0 = 1.15350369802766e-07 wbeta0 = 4.36024234050139e-06 pbeta0 = -5.46307999960091e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.52389060251324e-08 lagidl = -5.93862911325509e-15 wagidl = -4.60229080829501e-14 pagidl = 7.77807315977877e-21
+ bgidl = -2213402715.05922 lbgidl = 555.285556819766 wbgidl = 5461.95620038073 pbgidl = -0.000943842293977056
+ cgidl = -3324.35354454415 lcgidl = 0.000628238194704193 wcgidl = 0.00474696878500905 pcgidl = -8.22830075255898e-10
+ egidl = 19.278900492795 legidl = -3.32443225362009e-06 wegidl = -2.51194153250144e-05 pegidl = 4.35414921360734e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.967724069659923 lkt1 = 8.74187333149706e-08 wkt1 = 1.0054723644546e-06 pkt1 = -2.1394410814652e-13
+ kt2 = -0.398296571328263 lkt2 = 4.67586669004146e-08 wkt2 = 8.30760457021826e-07 pkt2 = -1.42063015348353e-13
+ at = -170851.234395878 lat = 0.0467967605966398 wat = 0.334981305312889 pat = -6.71413021064321e-8
+ ute = -0.942181992289765 lute = 6.2509323318015e-08 wute = 1.09154383237499e-06 pute = -1.06249734737074e-13
+ ua1 = -1.84132780195131e-09 lua1 = 3.33262721827451e-16 wua1 = 3.75631921824495e-15 pua1 = -6.35400242731618e-22
+ ub1 = 2.37210092666667e-19 wub1 = 2.64292757168557e-25
+ uc1 = 3.76355683135322e-12 luc1 = -7.46732450552953e-19 wuc1 = -5.37646616435935e-18 puc1 = 1.26925265831427e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.62 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.41151918892007 lvth0 = 3.62019446160894e-08 wvth0 = 9.57093991088551e-07 pvth0 = -1.29904219187719e-13
+ k1 = -2.26758269068731 lk1 = 5.19964047652529e-07 wk1 = 3.28050999080543e-06 pk1 = -4.78615118886645e-13
+ k2 = 1.270846046865 lk2 = -2.2836695526041e-07 wk2 = -1.52134750859296e-06 pk2 = 2.27252913095773e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 609409.86501181 lvsat = -0.0873951053415329 wvsat = -0.679172091022197 pvsat = 1.0784064138187e-7
+ ua = 1.51832618172493e-10 lua = -4.13271553606618e-16 wua = -1.68589330927599e-15 pua = 2.95482222769081e-22
+ ub = -1.92628253230173e-18 lub = 5.9226884219356e-25 wub = 3.72979820356283e-24 pub = -4.82201454889115e-31
+ uc = 2.58967002538763e-12 luc = -3.91639962880931e-19 wuc = -2.66739034501011e-18 puc = 4.39400747203288e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0106864132997624 lu0 = -1.29740353644785e-09 wu0 = -7.35355871177798e-09 pu0 = 1.34036116981227e-15
+ a0 = -0.855173815380581 la0 = 1.88491451404077e-07 wa0 = 3.63354841529781e-06 pa0 = -4.35779204973282e-13
+ keta = -0.832689077893654 lketa = 1.46599684637534e-07 wketa = 1.42392918628321e-06 pketa = -2.43627373490145e-13
+ a1 = 0.0
+ a2 = -3.2019090525702 la2 = 6.62794978372442e-07 wa2 = 3.92372605858992e-06 pa2 = -6.6537822287341e-13
+ ags = 1.25
+ b0 = 0.0
+ b1 = -4.08911049014536e-23 lb1 = 5.86124919436455e-30 wb1 = 6.95043366056275e-29 pb1 = -9.96261260037743e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.325624990069805 lvoff = -2.67320552947812e-08 wvoff = -3.46911122829019e-07 pvoff = 5.47018355928172e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -18.7383369998885 lnfactor = 3.44928078629959e-06 wnfactor = 2.51646927990893e-05 pnfactor = -3.74230710730038e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -2.40631671785476 leta0 = 4.31566335013593e-07 weta0 = 3.43301549625914e-06 peta0 = -5.66024376642542e-13
+ etab = -0.861273939966609 letab = 1.08466886342657e-07 wetab = 9.81422155772066e-07 petab = -1.23811849352912e-13
+ dsub = 0.37068240177151 ldsub = -1.58649941051246e-08 wdsub = -7.31692156842309e-08 pdsub = 1.04879290377462e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.71046415834999 lpclm = -5.28666775705477e-07 wpclm = -4.00898575898727e-06 ppclm = 6.86172022157109e-13
+ pdiblc1 = 3.47367782170907 lpdiblc1 = -5.54155971359683e-07 wpdiblc1 = -4.28707368099367e-06 ppdiblc1 = 7.14855098786177e-13
+ pdiblc2 = 0.0900650406287515 lpdiblc2 = -1.39171926141826e-08 wpdiblc2 = -1.17032870312573e-07 ppdiblc2 = 1.85924267276248e-14
+ pdiblcb = -0.986217486520106 lpdiblcb = 2.14462077171237e-07 wpdiblcb = 1.6746124030252e-06 ppdiblcb = -3.64292028791054e-13
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 9.62513689678327e-09 lpscbe2 = 2.59005612000915e-17 wpscbe2 = 1.00109926457981e-15 ppscbe2 = -2.6121158169936e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 15.8812623700667 lbeta0 = -1.3887199414252e-06 wbeta0 = -3.93890592882478e-06 pbeta0 = 8.92249762748357e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.21001594322295e-09 lagidl = -9.06819364237071e-16 wagidl = -9.88484558059839e-15 pagidl = 1.51397368174612e-21
+ bgidl = 942691899.894409 lbgidl = 8.21442845293495 wbgidl = 97.4089961512946 pbgidl = -1.39624106903343e-5
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.713698580275306 lkt1 = -2.04035705979502e-07 wkt1 = -1.32191798122296e-06 pkt1 = 1.89481079592537e-13
+ kt2 = -0.169356806016125 lkt2 = 7.07470586073925e-09 wkt2 = 6.46446916965319e-08 pkt2 = -9.26604081839745e-15
+ at = 573319.148647231 lat = -0.0821962452592865 wat = -0.622109915146003 pat = 9.87589758654713e-8
+ ute = -2.34524425071694 lute = 3.05713329069265e-07 wute = 2.76520966930472e-06 pute = -3.96359623578799e-13
+ ua1 = -2.37427591297519e-11 lua1 = 1.82061656748483e-17 wua1 = 2.46448790969746e-17 pua1 = 1.14407238676131e-23
+ ub1 = -3.92043284578177e-19 lub1 = 1.09073521904867e-25 wub1 = 1.52706593140277e-24 pub1 = -2.18886576475411e-31
+ uc1 = -3.3955526523995e-11 luc1 = 5.79141802009639e-18 wuc1 = 1.12435588772182e-17 puc1 = -1.61162924234271e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.63 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0053647
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29956891
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.7720538
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.64 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0053647
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29956891
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.7720538
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.65 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0074140810616 lvth0 = 1.63813955161699e-8
+ k1 = 0.533711539863405 lk1 = -3.35252744501912e-7
+ k2 = -0.015204835164966 lk2 = 1.01767887479373e-07 wk2 = 3.30872245021211e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67709.0584957215 lvsat = -0.0996868485549278
+ ua = -1.96104979334727e-09 lua = 4.53012753893265e-15
+ ub = 1.85327925148432e-18 lub = -2.29654397096517e-24
+ uc = -2.32886427786375e-11 luc = -1.24919512346539e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0046760248637794 lu0 = 2.0480533311125e-8
+ a0 = 1.3219165622399 la0 = -5.87602763891554e-7
+ keta = 0.0100523898791525 lketa = -2.72744888727377e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.199837851034395 lags = 4.15752045655893e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.318274014675695 lvoff = 1.49516223998211e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.4620747314211 lnfactor = 2.47776746807634e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0344627685079662 lpclm = 2.89382838858357e-07 wpclm = -9.92616735063633e-24 ppclm = -2.52435489670724e-29
+ pdiblc1 = 0.39
+ pdiblc2 = 9.85732448773808e-05 lpdiblc2 = 3.75099451691726e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799970624.466194 lpscbe1 = 0.117226568654587
+ pscbe2 = 1.20389481292726e-08 lpscbe2 = -1.01273764325456e-14
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.35955228517575e-10 lagidl = 8.59500572955045e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.629799548385 lkt1 = 6.72955516308661e-7
+ kt2 = -0.0781831266990001 lkt2 = 2.05421806009931e-7
+ at = -35193.10531325 lat = 0.361243766038403 wat = 1.38777878078145e-17 pat = -5.29395592033938e-23
+ ute = -2.44701888775 lute = 9.49223985116981e-6
+ ua1 = -2.428076454925e-09 lua1 = 1.73617415991573e-14 wua1 = 7.88860905221012e-31
+ ub1 = 2.00166536148e-18 lub1 = -1.20485610902818e-23
+ uc1 = 9.624331106095e-11 luc1 = -7.03799111305513e-16 wuc1 = -2.46519032881566e-32 puc1 = -2.82118644197349e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.66 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0087865031501 lvth0 = 2.18619407942096e-8
+ k1 = 0.438319171852289 lk1 = 4.56812235868604e-8
+ k2 = 0.01332183338898 lk2 = -1.21487420705046e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 32089.65415263 lvsat = 0.0425534723457048
+ ua = -6.30371477103069e-10 lua = -7.83720747101319e-16
+ ub = 1.12874327553622e-18 lub = 5.96773074155461e-25
+ uc = -6.4077122012637e-11 luc = 3.79626717408017e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104860229284 lu0 = -2.72075274025099e-9
+ a0 = 1.2151813426064 la0 = -1.61372955390757e-7
+ keta = 0.0112322389301054 lketa = -3.19860249221719e-08 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.231933635768609 lags = 2.87582728836931e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.28016803107749 lvoff = -2.65384833187796e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.3908807178428 lnfactor = -1.23126877212893e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.139268494014963 letab = 2.76612509352725e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.275233282675524 lpclm = 1.2508608823632e-06 ppclm = -2.01948391736579e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0018580315657347 lpdiblc2 = -3.27511725517847e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799999960.066619 lpscbe1 = 7.96007225289941e-5
+ pscbe2 = 9.63319118340849e-09 lpscbe2 = -5.20375801862541e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.038830824303e-12 lalpha0 = 1.21350786062605e-17
+ alpha1 = 2.9141211206745e-15 lalpha1 = -1.16370706077921e-20
+ beta0 = 56.9100629999999 lbeta0 = -0.000107460977160294
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.68775207909697e-11 lagidl = 3.6180069251305e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.451622277389999 lkt1 = -3.85665506919725e-8
+ kt2 = -0.00801757949699999 lkt2 = -7.4772939922609e-8
+ at = 102918.248221 lat = -0.190281550261352
+ ute = 0.75230175845 lute = -3.28372885948521e-06 wute = 4.2351647362715e-22 pute = -1.41363874215605e-27
+ ua1 = 3.98560513679e-09 lua1 = -8.25025682093871e-15
+ ub1 = -2.77182014511e-18 lub1 = 7.01357997563328e-24 pub1 = -2.80259692864963e-45
+ uc1 = -2.21393444354e-10 luc1 = 5.64631814289714e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.67 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.006776922084 lvth0 = 1.78561664910749e-8
+ k1 = 0.468810858652519 lk1 = -1.50990143961379e-8
+ k2 = 0.00448373627148799 lk2 = 5.46857276148265e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77900.294865342 lvsat = -0.0487626185912911
+ ua = -1.30087102961762e-09 lua = 5.52811489908928e-16
+ ub = 1.65098192376424e-18 lub = -4.44225068426082e-25
+ uc = -4.14092499588139e-11 luc = -7.22205900322166e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00867459456899998 lu0 = 8.90036242818672e-10
+ a0 = 1.6312399809578 la0 = -9.90718449444858e-7
+ keta = 0.0279922647790546 lketa = -6.53944213278645e-08 wketa = 6.61744490042422e-24 pketa = 2.52435489670724e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.393439099563341 lags = 1.53416196633805e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.2886710916924 lvoff = 1.42956255081255e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.4973376453944 lnfactor = 5.4986458881922e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.078470371 leta0 = 1.57414641388398e-07 weta0 = 2.31610571514848e-23 peta0 = 3.39210189245035e-29
+ etab = 0.00595669402992639 letab = -1.2870376534299e-08 petab = 4.73316543132607e-30
+ dsub = -0.0380014000000002 ldsub = 5.940175146732e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.333325541317719 lpclm = 3.77974532621591e-8
+ pdiblc1 = 0.39770896841646 lpdiblc1 = -1.536657968533e-8
+ pdiblc2 = 0.000215
+ pdiblcb = -0.4236676 lpdiblcb = 3.960116764488e-7
+ drout = 0.2110872461536 ldrout = 6.95501050926675e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.032799802395e-08 lpscbe2 = -1.90536067977383e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.32561383513941e-11 lalpha0 = 1.91968665957697e-16 walpha0 = 6.16297582203915e-33 palpha0 = -4.11423022787801e-38
+ alpha1 = -9.93396282422415e-11 lalpha1 = 1.98011627638892e-16 walpha1 = -4.42301848790681e-32 palpha1 = 5.21396029436995e-38
+ beta0 = -2.86171356345561 lbeta0 = 1.16843763911515e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9577639605148e-10 lagidl = -2.93805933700985e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.428378914775259 lkt1 = -8.48984286397128e-8
+ kt2 = -0.0273048137834199 lkt2 = -3.63269629045852e-8
+ at = -7927.86288261802 lat = 0.030672215153712 pat = -1.32348898008484e-23
+ ute = -0.598656317553001 lute = -5.90812790181536e-7
+ ua1 = -6.673817948866e-11 lua1 = -1.72566899554433e-16
+ ub1 = 1.01168299679436e-18 lub1 = -5.28220610244075e-25
+ uc1 = 7.6199295177312e-11 luc1 = -2.85711019421528e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.68 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.021883259604 lvth0 = 3.28618655905177e-8
+ k1 = 0.398846243563881 lk1 = 5.43994964267828e-8
+ k2 = 0.0243921037457624 lk2 = -1.43071651686781e-08 wk2 = 1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -12824.776391484 lvsat = 0.041358042240822
+ ua = -3.6513148601276e-10 lua = -3.76694156856437e-16
+ ub = 9.89933100099282e-19 lub = 2.12419847975621e-25
+ uc = -7.52043260124921e-11 luc = 2.63478742537868e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0117406951944 lu0 = -2.1556380202149e-9
+ a0 = 0.139135158719601 la0 = 4.9144597046759e-7
+ keta = -0.0422650138775481 lketa = 4.39480333832778e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.991513061907201 lags = 1.58436356167227e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.24715506755244 lvoff = -2.69438188790144e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.92532561224 lnfactor = 1.24727877808744e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32453716 leta0 = 4.0184213344008e-7
+ etab = -0.013900565275 letab = 6.85459370913795e-9
+ dsub = 0.799349363827521 ldsub = -2.37754818365702e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.11992164766228 lpclm = 2.49779650178066e-7
+ pdiblc1 = 0.60630129375168 lpdiblc1 = -2.22569262949166e-7
+ pdiblc2 = -9.79659804609995e-05 lpdiblc2 = 3.10881001099169e-10
+ pdiblcb = -0.025
+ drout = 0.823688067692801 ldrout = 8.69813760605692e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 7.5146551626052e-09 lpscbe2 = 8.89239691428671e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77191165332441 lbeta0 = 1.28254385565648e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.746561140738e-10 lagidl = 2.7282635504184e-16 pagidl = 9.4039548065783e-38
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.51916168720948 lkt1 = 5.27954896455041e-9
+ kt2 = -0.0724470689491601 lkt2 = 8.51455455724071e-9
+ at = -18539.604612764 lat = 0.0412132614604518 pat = 1.32348898008484e-23
+ ute = -2.133537872814 lute = 9.33843384158313e-7
+ ua1 = -1.02651999654268e-09 lua1 = 7.80820851034373e-16 wua1 = 3.94430452610506e-31
+ ub1 = 4.09283428091281e-19 lub1 = 7.01657725323038e-26
+ uc1 = 7.02451467413761e-11 luc1 = -2.2656620043097e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.69 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.948890704288003 lvth0 = -3.14813566396651e-9
+ k1 = 0.43987873475056 lk1 = 3.41566092897283e-8
+ k2 = 0.00505947892961119 lk2 = -4.76964670712773e-09 pk2 = 1.57772181044202e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 30780.1582495202 lvsat = 0.0198460709948983
+ ua = -7.20111477664003e-10 lua = -2.01569037735197e-16
+ ub = 1.1641954604768e-18 lub = 1.26449603631697e-25
+ uc = -4.30670652829792e-11 luc = 1.04933423200104e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00915178201416 lu0 = -8.78428769701665e-10
+ a0 = 1.44987763288 la0 = -1.55193100249753e-7
+ keta = -0.0561205618279248 lketa = 1.12302716530708e-8
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 2.17978636967648 lags = -4.27784020941055e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.18456167847128 lvoff = -5.78235162615357e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.356397574 lnfactor = 4.05401698337989e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 petab = 9.24446373305873e-33
+ dsub = 0.0151130540728808 ldsub = 1.49138754216033e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.615591804575359 lpclm = 5.24672630688115e-9
+ pdiblc1 = -0.14347143930832 lpdiblc1 = 1.47322117633188e-07 ppdiblc1 = -5.04870979341448e-29
+ pdiblc2 = -0.00972230637784599 lpdiblc2 = 5.05893384406429e-09 wpdiblc2 = 8.27180612553028e-25 ppdiblc2 = -1.97215226305253e-31
+ pdiblcb = 0.1696704 lpdiblcb = -9.60383057952e-08 wpdiblcb = -5.29395592033938e-23 ppdiblcb = 1.26217744835362e-29
+ drout = 1.55317580771432 ldrout = -2.72902646626167e-7
+ pscbe1 = 800069244.261281 lpscbe1 = -0.034160825371373
+ pscbe2 = 9.42176599694321e-09 lpscbe2 = -5.16105533619634e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77756825213281 lbeta0 = 1.2546377042271e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.493122281476e-10 lagidl = -1.33668538972981e-16
+ bgidl = 730034204.006401 lbgidl = 133.18438586389
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.504946199280001 lkt1 = -1.73349141960335e-9
+ kt2 = -0.0917821417920001 lkt2 = 1.80532807233817e-8
+ at = 63485.4642880001 lat = 0.000747178019086636
+ ute = -0.29451476672 lute = 2.65834030441113e-8
+ ua1 = 7.0578500184e-10 lua1 = -7.3791032257742e-17
+ ub1 = 6.6102183352e-19 lub1 = -5.40263489250896e-26
+ uc1 = 4.74348323563201e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.70 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.758071657257144 lvth0 = -4.95816609303614e-8
+ k1 = -0.777750412353429 lk1 = 3.30452050687719e-7
+ k2 = 0.462511999162372 lk2 = -1.16085228075527e-07 wk2 = -2.11758236813575e-22
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 237786.933100285 lvsat = -0.0305265435837374
+ ua = 1.09572681037143e-10 lua = -4.03462721545216e-16
+ ub = 3.70232301220002e-19 lub = 3.19651010878927e-25
+ uc = -3.747113248118e-13 luc = 1.04670292537848e-19 wuc = -1.92592994438724e-34 puc = 2.29588740394978e-41
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0106202771988571 lu0 = -1.2357694509555e-9
+ a0 = 0.131411673999997 la0 = 1.65639769252188e-7
+ keta = -0.101820143345726 lketa = 2.23507164204494e-08 wketa = 2.64697796016969e-23 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.119936524349429 la2 = 9.82566566797385e-8
+ ags = -1.62902379023886 lags = 4.99044225752423e-7
+ b0 = 0.0
+ b1 = -5.21832167044571e-24 lb1 = 1.26981595864292e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.220178493333428 lvoff = -4.91565917666102e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.873008799999994 lnfactor = 5.230285558256e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.17996084013057 leta0 = -1.67893690915693e-7
+ etab = 0.0779204436747429 letab = -1.89762135479246e-08 wetab = 2.35746474577613e-23 petab = 1.62702561701834e-30
+ dsub = 1.515770617532 ldsub = -2.16028255960982e-07 wdsub = -1.6940658945086e-21
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.674530623428858 lpclm = -9.09532799529139e-9
+ pdiblc1 = 1.228866610524 lpdiblc1 = -1.86619878736909e-07 ppdiblc1 = 2.01948391736579e-28
+ pdiblc2 = 0.03274100563686 lpdiblc2 = -5.27400357497024e-9
+ pdiblcb = -0.596438571428571 lpdiblcb = 9.03851190942857e-8
+ drout = -0.975627884694001 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066854 lpscbe1 = 0.0428666491488912
+ pscbe2 = 8.76724844606286e-09 lpscbe2 = 1.07658438434153e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.5332516765828 lbeta0 = -3.01760722716119e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1956850179.27428 lbgidl = -165.346559925846
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.20003683742857 lkt1 = -7.59295257138061e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080508e-08 wkt2 = 5.29395592033938e-23 pkt2 = 1.26217744835362e-29
+ at = 84910.017942857 lat = -0.00446623001817895
+ ute = -0.108778416857143 lute = -1.86133088588166e-8
+ ua1 = 1.02665585028571e-09 lua1 = -1.51871102776825e-16
+ ub1 = 4.39e-19
+ uc1 = -3.41423648285715e-13 luc1 = 2.22353418646549e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.71 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = 0.0887006526805187 lvth0 = -1.96359479590336e-07 wvth0 = -1.00780724473305e-06 pvth0 = 1.74691292187539e-13
+ k1 = 3.75173699010685 lk1 = -4.5468023667994e-07 wk1 = -4.60324701042119e-06 pk1 = 7.9791763029239e-13
+ k2 = -0.736579800550957 lk2 = 9.17629463031819e-08 wk2 = 1.10786283713848e-06 pk2 = -1.92034728463909e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -323162.505808177 lvsat = 0.0667073102577777 wvsat = 0.542257297594787 pvsat = -9.39937954504853e-8
+ ua = -1.31393747733486e-08 lua = 1.89308333230309e-15 wua = 1.57221619003511e-14 pua = -2.72524809948305e-21
+ ub = 1.03322383706342e-17 lub = -1.4071431971812e-24 wub = -1.23257039325945e-23 pub = 2.13651286826807e-30
+ uc = 1.91739534997083e-12 luc = -2.92638894255624e-19 wuc = -1.78688383262543e-18 puc = 3.09734869779627e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0253214631398974 lu0 = 4.99429993588354e-09 wu0 = 3.98074765936302e-08 pu0 = -6.90014837778667e-15
+ a0 = -1.68631396147731 la0 = 4.80720695454553e-07 wa0 = 4.72212773875486e-06 pa0 = -8.1852417798029e-13
+ keta = 0.642009079699266 lketa = -1.06583153443723e-07 wketa = -5.0754522297849e-07 pketa = 8.79768738606455e-14
+ a1 = 0.0
+ a2 = 2.22133314433735 la2 = -2.65995230635728e-07 wa2 = -3.17932310752062e-06 pa2 = 5.51097508811409e-13
+ ags = 1.25
+ b0 = 0.0
+ b1 = 1.21760838977067e-23 lb1 = -1.74529551372948e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.241123253568276 lvoff = -1.29117713971058e-07 wvoff = -1.08920521429769e-06 pvoff = 1.88800653435934e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -9.87283685517585 lnfactor = 2.38569195000247e-06 wnfactor = 1.3553173135453e-05 pnfactor = -2.34927992495316e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 2.75461061823134 leta0 = -4.40840334152124e-07 weta0 = -3.32646882694641e-06 peta0 = 5.76603453525237e-13
+ etab = 0.172175835684881 letab = -3.53142546881779e-08 wetab = -3.72130626979222e-07 petab = 6.45043786193245e-14
+ dsub = 0.43612777627507 ldsub = -2.88851251431879e-08 wdsub = -1.58885784466345e-07 pdsub = 2.75409441078276e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.48628077310331 lpclm = 5.38793397856802e-07 wpclm = 4.10715258037321e-06 ppclm = -7.11925613976732e-13
+ pdiblc1 = -2.16557451097412 lpdiblc1 = 4.01765756381333e-07 wpdiblc1 = 3.09889307556994e-06 ppdiblc1 = -5.37155927933143e-13
+ pdiblc2 = -0.0421335406898698 lpdiblc2 = 7.70460053621247e-09 wpdiblc2 = 5.6113190420557e-08 ppdiblc2 = -9.72654820111851e-15
+ pdiblcb = 3.22192240415097 lpdiblcb = -5.71481935690721e-07 wpdiblcb = -3.8369659952901e-06 ppdiblcb = 6.65092011691596e-13
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.41961622561841e-08 lpscbe2 = -8.33378623584643e-16 wpscbe2 = -4.98576554589766e-15 ppscbe2 = 8.64222628194804e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -0.376966146498177 lbeta0 = 1.5893946143011e-06 wbeta0 = 1.73551820565636e-05 pbeta0 = -3.00831254732062e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.67672932376725e-09 lagidl = -1.48667310752317e-15 wagidl = -1.31156041904019e-14 pagidl = 2.27343259915589e-21
+ bgidl = 1017064548.30667 lbgidl = -2.44599822518103
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.295597738666668 lkt1 = -5.93651902149972e-8
+ kt2 = -0.12
+ at = -477168.708323278 lat = 0.0929633722353404 wat = 0.753758361715837 pat = -1.306549669031e-7
+ ute = -0.233981691333334 lute = 3.08917633233733e-9
+ ua1 = -1.45964257110642e-09 lua1 = 2.79098892990444e-16 wua1 = 1.90530345781488e-15 pua1 = -3.30261490770716e-22
+ ub1 = 7.73885347333333e-19 lub1 = -5.80483563360657e-26
+ uc1 = 3.8082395871078e-12 luc1 = -4.96940907250094e-19 wuc1 = -3.82172392294229e-17 puc1 = 6.62449981354972e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0053647
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29956891
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.7720538
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0053647
+ k1 = 0.49177002
+ k2 = -0.002473247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.3943119e-9
+ ub = 1.565972e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0072382252
+ a0 = 1.248405
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.25185017
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.29956891
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.7720538
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0074140810616 lvth0 = 1.63813955161632e-8
+ k1 = 0.533711539863404 lk1 = -3.35252744501908e-7
+ k2 = -0.015204835164966 lk2 = 1.01767887479373e-07 wk2 = -3.30872245021211e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67709.0584957215 lvsat = -0.0996868485549274
+ ua = -1.96104979334726e-09 lua = 4.53012753893265e-15
+ ub = 1.85327925148432e-18 lub = -2.29654397096517e-24
+ uc = -2.32886427786375e-11 luc = -1.24919512346539e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00467602486377941 lu0 = 2.04805333111249e-8
+ a0 = 1.3219165622399 la0 = -5.87602763891561e-7
+ keta = 0.0100523898791525 lketa = -2.72744888727377e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.199837851034395 lags = 4.15752045655891e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.318274014675695 lvoff = 1.49516223998211e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.4620747314211 lnfactor = 2.47776746807634e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0344627685079662 lpclm = 2.89382838858357e-07 wpclm = 3.30872245021211e-24 ppclm = -2.52435489670724e-29
+ pdiblc1 = 0.39
+ pdiblc2 = 9.85732448773808e-05 lpdiblc2 = 3.75099451691725e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799970624.466194 lpscbe1 = 0.117226568647311
+ pscbe2 = 1.20389481292726e-08 lpscbe2 = -1.01273764325455e-14
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.35955228517575e-10 lagidl = 8.59500572955037e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.629799548385 lkt1 = 6.72955516308661e-7
+ kt2 = -0.078183126699 lkt2 = 2.05421806009932e-7
+ at = -35193.10531325 lat = 0.361243766038403 wat = 1.38777878078145e-17
+ ute = -2.44701888775 lute = 9.49223985116982e-6
+ ua1 = -2.428076454925e-09 lua1 = 1.73617415991573e-14 pua1 = -1.50463276905253e-36
+ ub1 = 2.00166536148e-18 lub1 = -1.20485610902818e-23 pub1 = 5.60519385729927e-45
+ uc1 = 9.624331106095e-11 luc1 = -7.03799111305513e-16 wuc1 = 1.23259516440783e-32 puc1 = 9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0087865031501 lvth0 = 2.1861940794213e-8
+ k1 = 0.43831917185229 lk1 = 4.56812235868587e-8
+ k2 = 0.01332183338898 lk2 = -1.21487420705046e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 32089.6541526299 lvsat = 0.0425534723457046
+ ua = -6.30371477103069e-10 lua = -7.83720747101323e-16
+ ub = 1.12874327553622e-18 lub = 5.96773074155464e-25
+ uc = -6.40771220126369e-11 luc = 3.79626717408019e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104860229284 lu0 = -2.72075274025099e-9
+ a0 = 1.2151813426064 la0 = -1.61372955390757e-7
+ keta = 0.0112322389301054 lketa = -3.19860249221718e-08 pketa = -1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.231933635768609 lags = 2.87582728836931e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.28016803107749 lvoff = -2.65384833187881e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.3908807178428 lnfactor = -1.23126877212893e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.139268494014963 letab = 2.76612509352725e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.275233282675524 lpclm = 1.2508608823632e-06 wpclm = 1.05879118406788e-22 ppclm = -8.07793566946316e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0018580315657347 lpdiblc2 = -3.27511725517847e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799999960.06662 lpscbe1 = 7.96007225289941e-5
+ pscbe2 = 9.63319118340849e-09 lpscbe2 = -5.20375801862541e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.038830824303e-12 lalpha0 = 1.21350786062605e-17
+ alpha1 = 2.9141211206745e-15 lalpha1 = -1.16370706077921e-20
+ beta0 = 56.910063 lbeta0 = -0.000107460977160294
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.68775207909697e-11 lagidl = 3.6180069251305e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.451622277389999 lkt1 = -3.85665506919708e-8
+ kt2 = -0.00801757949699999 lkt2 = -7.4772939922609e-8
+ at = 102918.248221 lat = -0.190281550261352
+ ute = 0.75230175845 lute = -3.28372885948521e-06 wute = 3.17637355220363e-22
+ ua1 = 3.98560513679e-09 lua1 = -8.2502568209387e-15
+ ub1 = -2.77182014511e-18 lub1 = 7.01357997563327e-24 wub1 = -1.46936793852786e-39 pub1 = -2.80259692864963e-45
+ uc1 = -2.21393444354e-10 luc1 = 5.64631814289713e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.006776922084 lvth0 = 1.78561664910766e-8
+ k1 = 0.46881085865252 lk1 = -1.50990143961371e-8
+ k2 = 0.00448373627148801 lk2 = 5.46857276148265e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77900.2948653419 lvsat = -0.0487626185912911
+ ua = -1.30087102961762e-09 lua = 5.52811489908926e-16
+ ub = 1.65098192376424e-18 lub = -4.44225068426085e-25
+ uc = -4.1409249958814e-11 luc = -7.22205900322166e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00867459456899999 lu0 = 8.90036242818685e-10
+ a0 = 1.6312399809578 la0 = -9.9071844944486e-7
+ keta = 0.0279922647790546 lketa = -6.53944213278646e-08 wketa = 6.61744490042422e-24
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.393439099563341 lags = 1.53416196633805e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.2886710916924 lvoff = 1.42956255081255e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.4973376453944 lnfactor = 5.49864588819217e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.0784703710000001 leta0 = 1.57414641388398e-07 weta0 = -1.24077091882954e-23 peta0 = -2.52435489670724e-29
+ etab = 0.00595669402992638 letab = -1.2870376534299e-08 wetab = 1.65436122510606e-24 petab = -5.52202633654708e-30
+ dsub = -0.0380014000000002 ldsub = 5.94017514673201e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.33332554131772 lpclm = 3.77974532621582e-8
+ pdiblc1 = 0.39770896841646 lpdiblc1 = -1.53665796853292e-8
+ pdiblc2 = 0.000215
+ pdiblcb = -0.423667599999999 lpdiblcb = 3.960116764488e-7
+ drout = 0.2110872461536 ldrout = 6.95501050926675e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.032799802395e-08 lpscbe2 = -1.90536067977383e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.32561383513941e-11 lalpha0 = 1.91968665957697e-16 walpha0 = -4.93038065763132e-32 palpha0 = -8.81620763116716e-38
+ alpha1 = -9.93396282422415e-11 lalpha1 = 1.98011627638891e-16 walpha1 = 1.17301170675335e-32 palpha1 = 4.12628363674874e-38
+ beta0 = -2.86171356345561 lbeta0 = 1.16843763911515e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9577639605148e-10 lagidl = -2.93805933700986e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.428378914775259 lkt1 = -8.48984286397136e-8
+ kt2 = -0.02730481378342 lkt2 = -3.63269629045852e-8
+ at = -7927.86288261801 lat = 0.030672215153712
+ ute = -0.598656317552999 lute = -5.90812790181536e-7
+ ua1 = -6.67381794886596e-11 lua1 = -1.72566899554434e-16
+ ub1 = 1.01168299679436e-18 lub1 = -5.28220610244075e-25
+ uc1 = 7.61992951773119e-11 luc1 = -2.85711019421528e-17 wuc1 = -9.86076131526265e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.77 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.021883259604 lvth0 = 3.28618655905177e-8
+ k1 = 0.39884624356388 lk1 = 5.43994964267828e-8
+ k2 = 0.0243921037457624 lk2 = -1.43071651686781e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -12824.776391484 lvsat = 0.041358042240822 pvsat = -2.64697796016969e-23
+ ua = -3.65131486012761e-10 lua = -3.76694156856437e-16
+ ub = 9.89933100099277e-19 lub = 2.12419847975622e-25
+ uc = -7.52043260124921e-11 luc = 2.63478742537868e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0117406951944 lu0 = -2.1556380202149e-09 wu0 = 1.32348898008484e-23
+ a0 = 0.139135158719601 la0 = 4.91445970467591e-7
+ keta = -0.0422650138775481 lketa = 4.39480333832778e-09 wketa = -5.29395592033938e-23
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.991513061907201 lags = 1.58436356167227e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.24715506755244 lvoff = -2.69438188790142e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.92532561224 lnfactor = 1.24727877808744e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.32453716 leta0 = 4.0184213344008e-07 weta0 = 1.05879118406788e-22 peta0 = -2.01948391736579e-28
+ etab = -0.013900565275 letab = 6.85459370913796e-9
+ dsub = 0.79934936382752 ldsub = -2.37754818365701e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.11992164766228 lpclm = 2.49779650178066e-7
+ pdiblc1 = 0.60630129375168 lpdiblc1 = -2.22569262949166e-7
+ pdiblc2 = -9.79659804609995e-05 lpdiblc2 = 3.10881001099169e-10 ppdiblc2 = -1.97215226305253e-31
+ pdiblcb = -0.025
+ drout = 0.8236880676928 ldrout = 8.69813760605692e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 7.51465516260521e-09 lpscbe2 = 8.89239691428677e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77191165332439 lbeta0 = 1.28254385565641e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.746561140738e-10 lagidl = 2.72826355041841e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.519161687209481 lkt1 = 5.27954896455041e-9
+ kt2 = -0.07244706894916 lkt2 = 8.51455455724071e-9
+ at = -18539.604612764 lat = 0.0412132614604517
+ ute = -2.133537872814 lute = 9.33843384158313e-7
+ ua1 = -1.02651999654268e-09 lua1 = 7.80820851034374e-16 pua1 = 1.88079096131566e-37
+ ub1 = 4.0928342809128e-19 lub1 = 7.01657725323045e-26
+ uc1 = 7.0245146741376e-11 luc1 = -2.2656620043097e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.78 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.948890704288001 lvth0 = -3.14813566396651e-9
+ k1 = 0.43987873475056 lk1 = 3.41566092897283e-8
+ k2 = 0.00505947892961119 lk2 = -4.76964670712773e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 30780.15824952 lvsat = 0.0198460709948983
+ ua = -7.20111477664003e-10 lua = -2.01569037735197e-16
+ ub = 1.1641954604768e-18 lub = 1.26449603631696e-25
+ uc = -4.30670652829792e-11 luc = 1.04933423200104e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00915178201416002 lu0 = -8.78428769701665e-10
+ a0 = 1.44987763288 la0 = -1.55193100249753e-7
+ keta = -0.0561205618279248 lketa = 1.12302716530708e-8
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 2.17978636967648 lags = -4.27784020941055e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.18456167847128 lvoff = -5.78235162615357e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.35639757400001 lnfactor = 4.05401698337989e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 wetab = -1.29246970711411e-26 petab = 9.24446373305873e-33
+ dsub = 0.0151130540728799 ldsub = 1.49138754216033e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.615591804575361 lpclm = 5.24672630688115e-9
+ pdiblc1 = -0.14347143930832 lpdiblc1 = 1.47322117633188e-7
+ pdiblc2 = -0.009722306377846 lpdiblc2 = 5.05893384406429e-09 ppdiblc2 = 1.57772181044202e-30
+ pdiblcb = 0.1696704 lpdiblcb = -9.60383057952e-08 wpdiblcb = -1.05879118406788e-22 ppdiblcb = 5.04870979341448e-29
+ drout = 1.55317580771432 ldrout = -2.72902646626167e-7
+ pscbe1 = 800069244.26128 lpscbe1 = -0.0341608253716004
+ pscbe2 = 9.42176599694321e-09 lpscbe2 = -5.16105533619603e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.77756825213281 lbeta0 = 1.2546377042271e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.493122281476e-10 lagidl = -1.33668538972981e-16
+ bgidl = 730034204.006401 lbgidl = 133.184385863891
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.50494619928 lkt1 = -1.73349141960335e-9
+ kt2 = -0.0917821417920001 lkt2 = 1.80532807233817e-8
+ at = 63485.464288 lat = 0.000747178019086692
+ ute = -0.29451476672 lute = 2.65834030441114e-8
+ ua1 = 7.0578500184e-10 lua1 = -7.3791032257742e-17
+ ub1 = 6.61021833520001e-19 lub1 = -5.402634892509e-26
+ uc1 = 4.74348323563201e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.79 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.75807165725714 lvth0 = -4.95816609303614e-8
+ k1 = -0.777750412353427 lk1 = 3.30452050687719e-7
+ k2 = 0.462511999162371 lk2 = -1.16085228075527e-07 wk2 = -5.29395592033938e-23 pk2 = -2.52435489670724e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 237786.933100285 lvsat = -0.0305265435837373
+ ua = 1.09572681037143e-10 lua = -4.03462721545216e-16
+ ub = 3.70232301220002e-19 lub = 3.19651010878929e-25
+ uc = -3.74711324811799e-13 luc = 1.04670292537848e-19 puc = 2.29588740394978e-41
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0106202771988571 lu0 = -1.2357694509555e-9
+ a0 = 0.131411673999999 la0 = 1.65639769252188e-7
+ keta = -0.101820143345726 lketa = 2.23507164204494e-08 pketa = -6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.119936524349429 la2 = 9.82566566797391e-8
+ ags = -1.62902379023885 lags = 4.99044225752423e-7
+ b0 = 0.0
+ b1 = -5.21832167044571e-24 lb1 = 1.26981595864292e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.22017849333343 lvoff = -4.91565917666104e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.873008800000008 lnfactor = 5.23028555825598e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.17996084013057 leta0 = -1.67893690915693e-7
+ etab = 0.0779204436747427 letab = -1.89762135479246e-08 wetab = -3.30872245021211e-24 petab = -4.95503256091948e-30
+ dsub = 1.515770617532 ldsub = -2.16028255960982e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.674530623428856 lpclm = -9.09532799529139e-9
+ pdiblc1 = 1.228866610524 lpdiblc1 = -1.86619878736909e-7
+ pdiblc2 = 0.0327410056368599 lpdiblc2 = -5.27400357497024e-9
+ pdiblcb = -0.596438571428571 lpdiblcb = 9.03851190942857e-08 ppdiblcb = -1.0097419586829e-28
+ drout = -0.975627884693997 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066856 lpscbe1 = 0.0428666491493459
+ pscbe2 = 8.76724844606284e-09 lpscbe2 = 1.07658438434153e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.5332516765829 lbeta0 = -3.01760722716119e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1956850179.27428 lbgidl = -165.346559925845
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.20003683742857 lkt1 = -7.59295257138064e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080507e-08 wkt2 = 5.29395592033938e-23
+ at = 84910.017942857 lat = -0.00446623001817897
+ ute = -0.108778416857143 lute = -1.86133088588166e-8
+ ua1 = 1.02665585028571e-09 lua1 = -1.51871102776825e-16
+ ub1 = 4.39e-19
+ uc1 = -3.41423648285712e-13 luc1 = 2.22353418646549e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.80 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.68809962941481 lvth0 = 1.11627527707503e-07 wvth0 = 8.57374992354309e-07 pvth0 = -1.48615666424711e-13
+ k1 = -4.79593045011757 lk1 = 1.02695534207368e-06 wk1 = 4.36960021314835e-06 pk1 = -7.57417761746708e-13
+ k2 = 0.774294181522594 lk2 = -1.70128928001483e-07 wk2 = -4.78165340726173e-07 pk2 = 8.28842238307933e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 201423.849894585 lvsat = -0.0242234394670275 wvsat = -0.00842313753061186 pvsat = 1.46004981328121e-9
+ ua = 8.19003938326279e-09 lua = -1.80411465877561e-15 wua = -6.66822424112128e-15 pua = 1.15585665350748e-21
+ ub = -5.11203448390804e-18 lub = 1.26993617087945e-24 wub = 3.88680103113297e-24 pub = -6.73730317134527e-31
+ uc = -1.84786167456466e-12 luc = 3.60023227863309e-19 wuc = 2.16566535987591e-18 puc = -3.7539210215017e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0302110942004943 lu0 = -4.63160248838528e-09 wu0 = -1.84873923204987e-08 pu0 = 3.2045676100506e-15
+ a0 = 11.3490942475238 la0 = -1.77881089267728e-06 wa0 = -8.96169035245999e-06 pa0 = 1.55340148231471e-12
+ keta = 2.73604915463084 lketa = -4.69559871952213e-07 wketa = -2.70574745812533e-06 pketa = 4.69008852896528e-13
+ a1 = 0.0
+ a2 = -0.807337235419329 la2 = 2.58988435650536e-7
+ ags = -16.580389915694 lags = 3.09068412720657e-06 wags = 1.87173127369585e-05 pags = -3.2444215551989e-12
+ b0 = 0.0
+ b1 = 1.21760838977067e-23 lb1 = -1.74529551372948e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -1.7617021702891 lvoff = 2.18048039349531e-07 wvoff = 1.01324515235828e-06 pvoff = -1.75633888219479e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 38.5196597012058 lnfactor = -6.00256661808762e-06 wnfactor = -3.72464726631354e-05 pnfactor = 6.45622907848257e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.16073378506698 leta0 = -1.6456091164508e-07 weta0 = -1.65330905357142e-06 peta0 = 2.86581284727963e-13
+ etab = -1.2852994633915 letab = 2.17321598703125e-07 wetab = 1.15784269991888e-06 petab = -2.00698137918539e-13
+ dsub = 0.11768710587126 ldsub = 2.63127437832675e-08 wdsub = 1.75394825452823e-07 pdsub = -3.04025882543413e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.04834640137308 lpclm = 6.36220729729829e-07 wpclm = 4.69717658953751e-06 ppclm = -8.14199195677253e-13
+ pdiblc1 = 0.786477026603333 lpdiblc1 = -1.09936953039269e-7
+ pdiblc2 = 0.01132071733706 lpdiblc2 = -1.5610536416595e-9
+ pdiblcb = -0.43322835123459 lpdiblcb = 6.20945859463013e-8
+ drout = 1.0
+ pscbe1 = -22426056.9391708 lpscbe1 = 142.557687857722 wpscbe1 = 863.33533834865 ppscbe1 = -0.000149648820878678
+ pscbe2 = -5.82203873378868e-09 lpscbe2 = 2.63653629961527e-15 wpscbe2 = 1.60281848013586e-14 ppscbe2 = -2.77829349709789e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.4098268772649 lbeta0 = -1.32039451485194e-06 wbeta0 = -2.66622983146096e-07 pbeta0 = 4.62158946525801e-14
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.23766860745942e-08 lagidl = 3.896063810798e-15 wagidl = 1.94824764073878e-14 pagidl = -3.37705349550379e-21
+ bgidl = 1017064548.30666 lbgidl = -2.44599822518103
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.295597738666672 lkt1 = -5.93651902149972e-8
+ kt2 = -0.12
+ at = 240872.694333334 lat = -0.0315004884183513
+ ute = -0.233981691333334 lute = 3.08917633233733e-9
+ ua1 = 3.55377781333335e-10 lua1 = -3.55131048607573e-17
+ ub1 = 7.73885347333335e-19 lub1 = -5.8048356336065e-26
+ uc1 = -3.25980697233334e-11 luc1 = 5.81365593600315e-18 wuc1 = -6.16297582203915e-33 puc1 = -2.93873587705572e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.81 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.965665208194601 wvth0 = -3.53223131778187e-8
+ k1 = 0.53696217035377 wk1 = -4.02093632784939e-8
+ k2 = 0.0032854709802425 wk2 = -5.12377440492052e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161274.634028667 wvsat = -0.0943454308640837
+ ua = -3.06755650285381e-09 wua = 1.48875633408128e-15
+ ub = 2.14389095287385e-18 wub = -5.14198880551676e-25
+ uc = 6.14166013797161e-11 wuc = -8.92706797696628e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0033077195627891 wu0 = 9.38317209432245e-9
+ a0 = 1.2396907970452 wa0 = 7.75339410825026e-9
+ keta = 0.0039938051129965 wketa = 2.3546423962153e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.31008900098943 wags = -5.18175456099637e-8
+ b0 = 7.3488582699e-08 wb0 = -6.53858932454902e-14
+ b1 = -7.7516677147e-09 wb1 = 6.89698588614615e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.13114231410195 wvoff = -1.49856249972842e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.738744457629098 wnfactor = 9.19378927561639e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00036344016320659 wpdiblc2 = 8.28597784255739e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 834086075.39378 wpscbe1 = -30.3409078179893
+ pscbe2 = 1.50971808672986e-08 wpscbe2 = -3.84832174279197e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.448711e-10 walpha0 = 3.0684637123042e-16
+ alpha1 = -3.448711e-10 walpha1 = 3.0684637123042e-16
+ beta0 = 123.115197 wbeta0 = -8.28485202322134e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.39325340101386e-09 wagidl = 3.14965299146862e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.61458422 wkt1 = 6.13692742460839e-8
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.82 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.9656652081946 wvth0 = -3.53223131778196e-8
+ k1 = 0.53696217035377 wk1 = -4.02093632784945e-8
+ k2 = 0.0032854709802425 wk2 = -5.12377440492052e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161274.634028667 wvsat = -0.0943454308640837
+ ua = -3.06755650285381e-09 wua = 1.48875633408128e-15
+ ub = 2.14389095287385e-18 wub = -5.14198880551675e-25
+ uc = 6.1416601379716e-11 wuc = -8.92706797696628e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0033077195627891 wu0 = 9.38317209432245e-9
+ a0 = 1.2396907970452 wa0 = 7.75339410825026e-9
+ keta = 0.0039938051129965 wketa = 2.35464239621531e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.31008900098943 wags = -5.18175456099636e-8
+ b0 = 7.34885826990001e-08 wb0 = -6.53858932454902e-14
+ b1 = -7.7516677147e-09 wb1 = 6.89698588614615e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.13114231410195 wvoff = -1.49856249972842e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.738744457629098 wnfactor = 9.19378927561638e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00036344016320659 wpdiblc2 = 8.28597784255739e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 834086075.393781 wpscbe1 = -30.3409078179893
+ pscbe2 = 1.50971808672986e-08 wpscbe2 = -3.84832174279196e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.448711e-10 walpha0 = 3.0684637123042e-16
+ alpha1 = -3.448711e-10 walpha1 = 3.0684637123042e-16
+ beta0 = 123.115197 wbeta0 = -8.28485202322134e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.39325340101386e-09 wagidl = 3.14965299146862e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.614584219999999 wkt1 = 6.13692742460839e-8
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.83 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.72515996207783 lvth0 = -1.92243972298452e-06 wvth0 = -2.5113340078368e-07 pvth0 = 1.72505096738126e-12
+ k1 = 0.667501357871833 lk1 = -1.04344384807726e-06 wk1 = -1.19038447012418e-07 pk1 = 6.3010751051556e-13
+ k2 = 0.0446385709964666 lk2 = -3.30549305777485e-07 wk2 = -5.32452038535666e-08 pk2 = 3.84650850626182e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 256146.501807898 lvsat = -0.7583429058507 wvsat = -0.167660745374951 pvsat = 5.86034089461667e-7
+ ua = -5.3916837571497e-09 lua = 1.8577534698599e-14 wua = 3.0523798103483e-15 pua = -1.24985709505373e-20
+ ub = 5.90316992781693e-19 lub = 1.24182417710151e-23 wub = 1.12371081857504e-24 pub = -1.30923658385982e-29
+ uc = 1.14852851320696e-10 luc = -4.27134007230733e-16 wuc = -1.22910316871228e-16 puc = 2.68892989550151e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0284101931192186 lu0 = 2.00652555772603e-07 wu0 = 2.94382043778722e-08 pu0 = -1.60306651643325e-13
+ a0 = 1.55649481432839 la0 = -2.53232158990239e-06 wa0 = -2.08714170085369e-07 pa0 = 1.7302984066363e-12
+ keta = 0.0303000374491662 lketa = -2.10274606569534e-07 wketa = -1.80151864937686e-08 pketa = 1.62822927319806e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.075526637590849 lags = 1.87493625272369e-06 wags = 1.10604932533931e-07 pags = -1.29829776660176e-12
+ b0 = 4.65955853583017e-07 lb0 = -3.13712355011351e-12 wb0 = -4.14580586269831e-13 pb0 = 2.7912312091498e-18
+ b1 = -1.65368460393553e-08 lb1 = 7.02228997392437e-14 wb1 = 1.47135297761173e-14 pb1 = -6.24802773043741e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.118207338180848 lvoff = -1.99313605087888e-06 wvoff = -3.88355879149557e-07 pvoff = 1.90640814888414e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -1.9804230014034 lnfactor = 2.17352245786479e-05 wnfactor = 3.06293550629829e-06 pnfactor = -1.71341722559656e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.21129242978291 lpclm = -9.6683595263376e-06 wpclm = -1.10840097078876e-06 ppclm = 8.85982359904266e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00385536529229361 lpdiblc2 = 2.79121378274862e-08 wpdiblc2 = 3.5179859727273e-09 ppdiblc2 = -2.14971888036609e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 868115469.255025 lpscbe1 = -272.008447068059 wpscbe1 = -60.6313441210723 ppscbe1 = 0.000242121695538007
+ pscbe2 = 2.09454004135187e-08 lpscbe2 = -4.67467955311434e-14 wpscbe2 = -7.92444644958011e-15 ppscbe2 = 3.25818425115085e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.15893687774676e-10 lalpha0 = 2.16637514971765e-15 walpha0 = 5.47986604726753e-16 palpha0 = -1.92751539173511e-21
+ alpha1 = -6.89167701418303e-10 lalpha1 = 2.75207910738777e-15 walpha1 = 6.13181586828864e-16 palpha1 = -2.44864091958123e-21
+ beta0 = 194.26704357092 lbeta0 = -0.000568740758965504 wbeta0 = -0.000146155320734286 pbeta0 = 5.06032654111637e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.13596854634974e-09 lagidl = 2.99167871943888e-14 wagidl = 6.47013745768275e-15 pagidl = -2.65417546621991e-20
+ bgidl = 2107368073.11315 lbgidl = -8851.56729880212 wbgidl = -985.272105581455 pbgidl = 0.00787561296188425
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.532375164970481 lkt1 = -6.57124763511551e-07 wkt1 = -8.66825852328784e-08 pkt1 = 1.18342855434385e-12
+ kt2 = -0.187620131271737 lkt2 = 1.08018877326737e-06 wkt2 = 9.73707212099572e-08 pkt2 = -7.78317085934957e-13
+ at = -9258.91033287105 lat = 0.153942979802331 wat = -0.0230747476970713 pat = 1.84444257607413e-7
+ ute = -3.4587347911921 lute = 1.75792270273579e-05 wute = 9.00166333703561e-07 pute = -7.19533376151336e-12
+ ua1 = -7.74708200901268e-09 lua1 = 5.98783508168574e-14 wua1 = 4.73254370350619e-15 pua1 = -3.78288214218968e-20
+ ub1 = 6.95549342879971e-18 lub1 = -5.1646183226255e-23 wub1 = -4.40762988303878e-24 pub1 = 3.52316754340295e-29
+ uc1 = 2.18816134008649e-10 luc1 = -1.68356511474062e-15 wuc1 = -1.09058213149696e-16 puc1 = 8.71739159381564e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.84 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.48369657877072 lvth0 = 1.10665337284664e-06 wvth0 = 4.22547535484859e-07 pvth0 = -9.65184715295479e-13
+ k1 = 0.310784755338068 lk1 = 3.81046116051721e-07 wk1 = 1.1347275232508e-07 pk1 = -2.98388297224449e-13
+ k2 = -0.0809058222230736 lk2 = 1.70791890353048e-07 wk2 = 8.38383216051109e-08 pk2 = -1.62770000761923e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6328.02789852174 lvsat = 0.23926669911362 wvsat = 0.022921206018908 pvsat = -1.75024059153584e-7
+ ua = 9.28935636043634e-10 lua = -6.66283490777689e-15 wua = -1.3873813413268e-15 pua = 5.23089596737064e-21
+ ub = 5.29866001719286e-18 lub = -6.38376334540092e-24 wub = -3.71015089553841e-24 pub = 6.21087783111622e-30
+ uc = -1.28738524394411e-11 luc = 8.29218925093662e-17 wuc = -4.55577097172483e-17 puc = -4.00021159969081e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0423301789367373 lu0 = -8.1837660092584e-08 wu0 = -2.83330894240013e-08 pu0 = 7.0393651204861e-14
+ a0 = 0.805977799876988 la0 = 4.6474652355295e-07 wa0 = 3.64085660355861e-07 pa0 = -5.57084922658227e-13
+ keta = -0.0415269255683224 lketa = 7.65547342727979e-08 wketa = 4.6942055090993e-08 pketa = -9.65732938758026e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = 1.38197925172107 lags = -3.34217061648187e-06 wags = -1.0232441164379e-06 pags = 3.22954472692131e-12
+ b0 = -7.0518677536023e-07 lb0 = 1.53964481346546e-12 wb0 = 6.27434432919917e-13 pb0 = -1.36988696355135e-18
+ b1 = 3.32697706660904e-09 lb1 = -9.10005989508186e-15 wb1 = -2.96015189459428e-15 pb1 = 8.09670731118191e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.564367221686601 lvoff = 7.32614876873084e-07 wvoff = 2.5286401309077e-07 pvoff = -6.54199613155058e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 6.67145586754464 lnfactor = -1.28146520801193e-05 wnfactor = -3.80860835096105e-06 pnfactor = 1.03062249478946e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.1392684888935 letab = 2.76612488900993e-07 wetab = -4.55678155815718e-15 petab = 1.81967689549841e-20
+ dsub = 0.859000699999999 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.94416912670563 lpclm = 6.92580301472722e-06 wpclm = 2.3746648495262e-06 ppclm = -5.04923549772225e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00629790356823405 lpdiblc2 = -1.26332965374756e-08 wpdiblc2 = -3.95034148322218e-09 ppdiblc2 = 8.3263670226255e-15
+ pdiblcb = 0.462444668731799 lpdiblcb = -2.74519891854411e-06 wpdiblcb = -6.11648531935703e-07 ppdiblcb = 2.44251932522306e-12
+ drout = 0.56
+ pscbe1 = 799999822.347933 lpscbe1 = 0.000354120616975706 wpscbe1 = 0.000122534127513063 ppscbe1 = -2.44251931180717e-10
+ pscbe2 = 9.64315525817299e-09 lpscbe2 = -1.61311046698578e-15 wpscbe2 = -8.86545780193426e-18 ppscbe2 = 9.72252144963023e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.47298006479066e-10 lalpha0 = 2.95114208964001e-16 walpha0 = 1.28353476317255e-16 palpha0 = -2.51778473998583e-22
+ alpha1 = 1.09856605183185e-14 lalpha1 = -4.43325141949713e-20 walpha1 = -7.18158922104643e-21 palpha1 = 2.90905159072328e-26
+ beta0 = 100.526597136953 lbeta0 = -0.00019440347208378 wbeta0 = -3.88074710393879e-05 pbeta0 = 7.73564067067115e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.18678047687567e-10 lagidl = -1.84880532615097e-15 wagidl = -6.68908654762138e-16 pagidl = 1.96686946237936e-21
+ bgidl = -1214736146.2263 lbgidl = 4414.71772024643 wbgidl = 1970.54421116291 pbgidl = -0.00392796065679104
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.990108369035007 lkt1 = 1.17075863414108e-06 wkt1 = 4.7911379984963e-07 pkt1 = -1.07598765046876e-12
+ kt2 = 0.169707816943784 lkt2 = -3.46742500803708e-07 wkt2 = -1.58129785225095e-07 pkt2 = 2.41982795431383e-13
+ at = 162669.829780976 lat = -0.532626591386421 wat = -0.0531635036306529 pat = 3.0459883004971e-7
+ ute = 2.53384282221434 lute = -6.35116087420737e-06 wute = -1.58511226546402e-06 pute = 2.72922370912933e-12
+ ua1 = 1.51200806020696e-08 lua1 = -3.14379585901566e-14 wua1 = -9.90681269632386e-15 pua1 = 2.06310767850878e-20
+ ub1 = -1.34715955358992e-17 lub1 = 2.9926087365858e-23 wub1 = 9.52004169570669e-24 pub1 = -2.03862247328948e-29
+ uc1 = -5.20614354072123e-10 luc1 = 1.26923075167087e-15 wuc1 = 2.66229470498604e-16 puc1 = -6.26911408663171e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.85 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.859423135614458 lvth0 = -1.37734603787577e-07 wvth0 = -1.3110688215174e-07 pvth0 = 1.38435674247424e-13
+ k1 = 0.657368028317915 lk1 = -3.09811492143383e-07 wk1 = -1.67767270963862e-07 pk1 = 2.62218128318286e-13
+ k2 = -0.0455948556104336 lk2 = 1.00405198787341e-07 wk2 = 4.4557036513923e-08 pk2 = -8.44691225008245e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 762849.569148904 lvsat = -1.26873643687933 wvsat = -0.60942827418946 pvsat = 1.085462189026e-6
+ ua = -4.96352633601228e-09 lua = 5.0828334546771e-15 wua = 3.25881899015326e-15 pua = -4.03055170898115e-21
+ ub = 3.13693157806079e-18 lub = -2.07470790199829e-24 wub = -1.32211211450305e-24 pub = 1.45070938340477e-30
+ uc = 1.86582307318966e-10 luc = -3.14661650071138e-16 wuc = -2.02853709753758e-16 puc = 2.73541978123868e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0099876454102004 lu0 = 2.24494472554921e-08 wu0 = 1.66045824560217e-08 pu0 = -1.91823177851203e-14
+ a0 = 3.45437665409091 la0 = -4.81440755170812e-06 wa0 = -1.62212163445413e-06 pa0 = 3.40209755396374e-12
+ keta = 0.163032746319274 lketa = -3.3120183296828e-07 wketa = -1.20151215134654e-07 pketa = 2.36500071209249e-13
+ a1 = 0.0
+ a2 = -0.570294274927202 la2 = 2.73145964939484e-06 wa2 = 1.21920864282113e-06 pa2 = -2.43029491766379e-12
+ ags = -4.12625971097633 lags = 7.63761142094344e-06 wags = 3.32124802300394e-06 pags = -5.4304965453294e-12
+ b0 = 5.57355890638085e-07 lb0 = -9.77029459290286e-13 wb0 = -4.95903056319289e-13 pb0 = 8.6930434057375e-19
+ b1 = -9.72774657807711e-09 lb1 = 1.69224168253695e-14 wb1 = 8.6551866414208e-15 pb1 = -1.50565883755213e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.0691986110760774 lvoff = -2.54423531064076e-07 wvoff = -1.95273927743024e-07 pvoff = 2.39090773550695e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 7.84014345782272 lnfactor = -1.5144241463949e-05 wnfactor = -5.64346199772277e-06 pnfactor = 1.39637084464233e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.32608126080038 leta0 = -2.64233149924131e-06 weta0 = -1.24968885889166e-06 peta0 = 2.49105229060539e-12
+ etab = -0.535309554809244 letab = 1.06605619515135e-06 wetab = 4.81587423027911e-07 petab = -9.59966501530046e-13
+ dsub = -1.0657221061954 ldsub = 2.64261225171933e-06 wdsub = 9.1440648211585e-07 pdsub = -1.82272118824784e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.73893377609808 lpclm = -2.40920395934172e-06 wpclm = -1.25062896315159e-06 ppclm = 2.17720042025328e-12
+ pdiblc1 = 0.426036787903175 lpdiblc1 = -7.18334987253389e-08 wpdiblc1 = -2.52044564313128e-08 ppdiblc1 = 5.02410007738801e-14
+ pdiblc2 = 0.00044351946819426 lpdiblc2 = -9.6353024427052e-10 wpdiblc2 = -2.03323414373991e-10 ppdiblc2 = 8.5729351930379e-16
+ pdiblcb = -2.4837040749272 lpdiblcb = 3.12747132584364e-06 wpdiblcb = 1.83290138528197e-06 ppdiblcb = -2.43029491766379e-12
+ drout = 0.132697301170835 ldrout = 8.51758707078729e-07 wdrout = 6.97468421068433e-08 pdrout = -1.39029030751571e-13
+ pscbe1 = 795876407.695818 lpscbe1 = 8.21971323643265 wpscbe1 = 3.66893408862597 ppscbe1 = -7.31342573835267e-6
+ pscbe2 = 1.13026784410869e-08 lpscbe2 = -4.92110108936893e-15 wpscbe2 = -8.67214298640282e-16 ppscbe2 = 2.68323150666203e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.78343046749665e-11 lalpha0 = 1.96516332537222e-16 walpha0 = 4.0733877767013e-18 palpha0 = -4.04625086733295e-24
+ alpha1 = -9.93562343796287e-11 lalpha1 = 1.98028123146192e-16 walpha1 = 1.47751812125238e-20 palpha1 = -1.4676748955295e-26
+ beta0 = -6.20685847615589 lbeta0 = 1.83523808611436e-05 wbeta0 = 2.97631659394476e-06 pbeta0 = -5.93280496674065e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.49936455062403e-09 lagidl = -3.20564359854133e-15 wagidl = -9.81908952543322e-16 pagidl = 2.59078484995791e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.308869546253552 lkt1 = -1.87180598384462e-07 wkt1 = -1.06332528469114e-07 pkt1 = 9.10047627294653e-14
+ kt2 = 0.0692276212061779 lkt2 = -1.464515083925e-07 wkt2 = -8.58889810790018e-08 pkt2 = 9.79824553764174e-14
+ at = -60385.6255734575 lat = -0.0880016761211245 wat = 0.0466738851836254 pat = 1.05589169105434e-7
+ ute = 3.35565372383641 lute = -7.98930777322491e-06 wute = -3.5183165157079e-06 pute = 6.58275320290197e-12
+ ua1 = 3.20082681823455e-09 lua1 = -7.67885709119445e-15 wua1 = -2.90729046971724e-15 pua1 = 6.67866314894821e-21
+ ub1 = -7.15013116341382e-19 lub1 = 4.49790687882139e-24 wub1 = 1.53631439843284e-24 pub1 = -4.47195772960159e-30
+ uc1 = 1.29507157777217e-11 luc1 = 2.0565522246652e-16 wuc1 = 5.62749301818661e-17 puc1 = -2.08401045177286e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.86 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.02429016494824 lvth0 = 2.6034081396777e-08 wvth0 = 2.14152525617169e-09 pvth0 = 6.07496772966427e-15
+ k1 = 0.277808267571465 lk1 = 6.72196414769748e-08 wk1 = 1.07692595043038e-07 pk1 = -1.14066240612767e-14
+ k2 = 0.0902011196598536 lk2 = -3.44861036956955e-08 wk2 = -5.85530585992385e-08 pk2 = 1.79540531586932e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1028975.22170011 lvsat = 0.511151217213039 wvsat = 0.904111932739872 pvsat = -4.17994813044765e-7
+ ua = -8.66142550562498e-10 lua = 1.01274644000598e-15 wua = 4.45770686796826e-16 pua = -1.23624393342168e-21
+ ub = 2.1933894081532e-18 lub = -1.13745161002662e-24 wub = -1.07076586313177e-24 pub = 1.20103760076012e-30
+ uc = -2.07502846058195e-10 luc = 7.67981080142249e-17 wuc = 1.17711576282208e-16 puc = -4.48877019765265e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011010498421116 lu0 = 1.59119305837996e-09 wu0 = 6.49686883494607e-10 pu0 = -3.33371372689737e-15
+ a0 = -3.99208702022471 la0 = 2.58244778160921e-06 wa0 = 3.67572271018271e-06 pa0 = -1.86045255164913e-12
+ keta = -0.223389161120479 lketa = 5.26457317241094e-08 wketa = 1.61153797241049e-07 pketa = -4.29308871740078e-14
+ a1 = 0.0
+ a2 = 3.5405885498544 la2 = -1.35203647400807e-06 wa2 = -2.43841728564227e-06 pa2 = 1.20296390686419e-12
+ ags = 4.15204655216979 lags = -5.85544765877597e-07 wags = -2.81206002079992e-06 pags = 6.6195140028663e-13
+ b0 = -7.63776618893518e-07 lb0 = 3.35301665462817e-13 wb0 = 6.7956428920288e-13 pb0 = -2.98332041492551e-19
+ b1 = 7.07121378167302e-08 lb1 = -6.29815770595996e-14 wb1 = -6.29155730677607e-14 pb1 = 5.60373669324776e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.502899797474587 lvoff = 1.76388338030647e-07 wvoff = 2.27546878639337e-07 pvoff = -1.80913200619547e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -16.2897037903437 lnfactor = 8.82485274185011e-06 wnfactor = 1.62066803337195e-05 pnfactor = -7.74086823680687e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -3.13364042360076 leta0 = 1.78767951929836e-06 weta0 = 2.49937771778332e-06 peta0 = -1.23303800453579e-12
+ etab = 1.06863191191749 letab = -5.27199813524051e-07 wetab = -9.63174827828696e-07 petab = 4.75170743211353e-13
+ dsub = 2.78751565154149 ldsub = -1.18495523607552e-06 wdsub = -1.76895544679646e-06 pdsub = 8.42764183494051e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.96633750457257 lpclm = 1.27138280405711e-06 wpclm = 1.85623280787957e-06 ppclm = -9.08963437659276e-13
+ pdiblc1 = 0.689231955458777 lpdiblc1 = -3.33275260074686e-07 wpdiblc1 = -7.37869093947287e-08 ppdiblc1 = 9.84997974356532e-14
+ pdiblc2 = -0.000195366777709762 lpdiblc2 = -3.2890025853671e-10 wpdiblc2 = 8.66615996258679e-11 ppdiblc2 = 5.69240385467198e-16
+ pdiblcb = 0.6647422 wpdiblcb = -6.1369274246084e-7
+ drout = 0.420328173142241 ldrout = 5.66044031976397e-07 wdrout = 3.58886319969184e-07 pdrout = -4.26242261412392e-13
+ pscbe1 = 808247184.608363 lpscbe1 = -4.06864956032086 wpscbe1 = -7.33786817725104 ppscbe1 = 3.62004921082874e-6
+ pscbe2 = -2.48817233168534e-08 lpscbe2 = 3.102224018406e-14 wpscbe2 = 2.88244250603462e-14 ppscbe2 = -2.68106021509148e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 15.5543404033212 lbeta0 = -3.26384491139844e-06 wbeta0 = -6.03461307736544e-06 pbeta0 = 3.01809389109928e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.97571285711779e-09 lagidl = 2.23295884351012e-15 wagidl = 3.3819605888808e-15 pagidl = -1.74401259258124e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.489498227233902 lkt1 = -7.75526567680261e-09 wkt1 = -2.63928321382829e-08 pkt1 = 1.15976246555895e-14
+ kt2 = -0.170374632876666 lkt2 = 9.15545154736435e-08 wkt2 = 8.71302861694994e-08 pkt2 = -7.38841575136742e-14
+ at = -357041.480976851 lat = 0.206677857973572 wat = 0.301179404180311 pat = -1.47220834123696e-7
+ ute = -8.56891076383874 lute = 3.85581526583335e-06 wute = 5.72582283388071e-06 pute = -2.59980169033969e-12
+ ua1 = -1.03770323445347e-08 lua1 = 5.80854637383246e-15 wua1 = 8.31954542762961e-15 pua1 = -4.47337956765052e-21
+ ub1 = 6.77754494824054e-18 lub1 = -2.94473576393429e-24 wub1 = -5.66611101511295e-24 pub1 = 2.68248512583916e-30
+ uc1 = 4.13043360831461e-10 luc1 = -1.91772005385871e-16 wuc1 = -3.05002037160583e-16 puc1 = 1.50469095008728e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.87 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.980951512537821 lvth0 = 4.65347729392831e-09 wvth0 = 2.85258540659735e-08 pvth0 = -6.94142427670586e-15
+ k1 = 0.252308782950744 lk1 = 7.97995062207916e-08 wk1 = 1.66888901568262e-07 pk1 = -4.06104115298177e-14
+ k2 = 0.0542080779936456 lk2 = -1.67293685061717e-08 wk2 = -4.37295826581519e-08 pk2 = 1.06410691848694e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -95269.655412271 lvsat = 0.0505187805517312 wvsat = 0.112151838517032 pvsat = -2.72908040810576e-8
+ ua = 3.84897972353431e-09 lua = -1.31340255245239e-15 wua = -4.06531325735483e-15 pua = 9.89245197418209e-22
+ ub = -1.86044745912135e-18 lub = 8.62460162400871e-25 wub = 2.69115244549768e-24 pub = -6.54859653782514e-31
+ uc = -1.02337679370456e-10 luc = 2.49161350108288e-17 wuc = 5.27355665735425e-17 puc = -1.28325672988727e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0226981710655859 lu0 = -4.17477998869755e-09 wu0 = -1.20527939966716e-08 pu0 = 2.93290278556207e-15
+ a0 = 1.66152932818236 la0 = -2.06696000481239e-07 wa0 = -1.8831544501205e-07 pa0 = 4.58243037583423e-14
+ keta = -0.22053854649493 lketa = 5.12394152059706e-08 wketa = 1.46289619397188e-07 pketa = -3.55978234048729e-14
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 5.44070696557385 lags = -1.22128991690553e-06 wags = -2.90137866501904e-06 pags = 7.06015681588403e-13
+ b0 = -1.65993456595493e-07 lb0 = 4.03925157410342e-14 wb0 = 1.47691383256879e-13 pb0 = -3.59389258189624e-20
+ b1 = -1.12386369653478e-07 lb1 = 2.7347874418738e-14 wb1 = 9.99948957854986e-14 pb1 = -2.43325579506517e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.124092574886034 lvoff = -1.32930824964998e-07 wvoff = -2.74622714421495e-07 pvoff = 6.68261420818977e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 0.21223232851807 lnfactor = 6.83820580843069e-07 wnfactor = 1.01801210267863e-06 pnfactor = -2.47721029041613e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 wetab = -6.46234853557053e-27 petab = -3.08148791101958e-33
+ dsub = 0.14966330342655 ldsub = 1.16397565638811e-07 wdsub = -1.19715034870482e-07 pdsub = 2.91312171553135e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.585080749510564 lpclm = 1.26712254242382e-08 wpclm = 2.71469732576727e-08 ppclm = -6.60589017857557e-15
+ pdiblc1 = -0.422644040669374 lpdiblc1 = 2.15255420103184e-07 wpdiblc1 = 2.48391644514707e-07 ppdiblc1 = -6.04431259929198e-14
+ pdiblc2 = -0.0124736374744419 lpdiblc2 = 5.72843725044776e-09 wpdiblc2 = 2.44797538281369e-09 ppdiblc2 = -5.95685433703119e-16
+ pdiblcb = 1.5307745498544 lpdiblcb = -4.2724666741247e-07 wpdiblcb = -1.21103180072058e-06 ppdiblcb = 2.94690056323745e-13
+ drout = 2.67345537674649 ldrout = -5.45509236395318e-07 wdrout = -9.96760008365738e-07 pdrout = 2.42549586915702e-13
+ pscbe1 = 800069244.26128 lpscbe1 = -0.0341608253711456
+ pscbe2 = 6.60243097022716e-08 lpscbe2 = -1.38251603335292e-14 wpscbe2 = -5.0361671761975e-14 ppscbe2 = 1.22549084832155e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.59329040294026 lbeta0 = 1.70305573689528e-07 wbeta0 = 1.63959778951856e-07 pbeta0 = -3.98976446905875e-14
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.89019256021353e-10 lagidl = -2.16332167721724e-16 wagidl = -3.02251678335855e-16 pagidl = 7.35493189028902e-23
+ bgidl = 730034204.006402 lbgidl = 133.184385863891
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.498549009775686 lkt1 = -3.29017071920441e-09 wkt1 = -5.6918494633865e-09 pkt1 = 1.38504326472157e-15
+ kt2 = 0.0471321477421401 lkt2 = -1.57498446632769e-08 wkt2 = -1.23597905581543e-07 pkt2 = 3.00760671484015e-14
+ at = 57360.4956136553 lat = 0.0022376156463644 wat = 0.00544964310324264 pat = -1.32610525345685e-9
+ ute = -1.30588320526931 lute = 2.72687776143824e-07 wute = 8.9985717952543e-07 pute = -2.18969446351359e-13
+ ua1 = 2.36483485009753e-09 lua1 = -4.77500904233033e-16 wua1 = -1.47612666189832e-15 pua1 = 3.59197709653013e-22
+ ub1 = 1.16823729496324e-18 lub1 = -1.77451144881766e-25 wub1 = -4.51291000538526e-25 pub1 = 1.09816249489044e-31
+ uc1 = 4.743483235632e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.88 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.708437786079259 lvth0 = -6.16594678750467e-08 wvth0 = -4.41613497363315e-08 pvth0 = 1.07461345221392e-14
+ k1 = -2.02711795768269 lk1 = 6.34470650433051e-07 wk1 = 1.11161502838986e-06 pk1 = -2.70498177778332e-13
+ k2 = 0.545014304567405 lk2 = -1.36161174068177e-07 wk2 = -7.34057827161471e-08 pk2 = 1.78624163545817e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 738412.672293368 lvsat = -0.152347809707504 wvsat = -0.445427846566279 pvsat = 1.08389521327745e-7
+ ua = 5.86452439728656e-09 lua = -1.80386116227392e-15 wua = -5.12042340090954e-15 pua = 1.24599358953053e-21
+ ub = 1.32705326660253e-18 lub = 8.68201108046759e-26 wub = -8.51323990745568e-25 pub = 2.07159477260045e-31
+ uc = -1.68800651054782e-12 luc = 4.2424491644448e-19 wuc = 1.16849414780618e-18 puc = -2.8433902893886e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0375241069894086 lu0 = -7.78249358452872e-09 wu0 = -2.39374727062708e-08 pu0 = 5.82489673339853e-15
+ a0 = 1.95638728836938 la0 = -2.78446146797227e-07 wa0 = -1.62375781807536e-06 pa0 = 3.95121979934823e-13
+ keta = 0.182152680668966 lketa = -4.67506626296377e-08 wketa = -2.52662605179045e-07 pketa = 6.14824130190584e-14
+ a1 = 0.0
+ a2 = -0.0353204792273516 la2 = 1.36036585416105e-07 wa2 = 1.38138707927813e-07 pa2 = -3.36143969097381e-14
+ ags = -1.62902379023885 lags = 4.99044225752423e-7
+ b0 = -4.26994762369998e-09 lb0 = 1.0390405148559e-15 wb0 = 3.79915259259559e-15 pb0 = -9.24478193577026e-22
+ b1 = 6.44215537882842e-10 lb1 = -1.56762120557335e-16 wb1 = -5.73185749950068e-16 pb1 = 1.3947787402135e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.412683937009636 lvoff = -2.03156069841431e-07 wvoff = -5.63084411070787e-07 pvoff = 1.37019834421143e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 23.1890864511252 lnfactor = -4.90732114764391e-06 wnfactor = -1.9855556024683e-05 pnfactor = 4.83161129193432e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.430993751557764 leta0 = 1.43584624834372e-08 weta0 = 6.66387625114366e-07 peta0 = -1.62157431920079e-13
+ etab = -0.497100985801246 letab = 1.20948351057903e-07 wetab = 5.11620831709111e-07 petab = -1.24496789946432e-13
+ dsub = 1.44415360420511 ldsub = -1.98601115172043e-07 wdsub = 6.37206789948942e-08 pdsub = -1.55056625852597e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.708064400894729 lpclm = -1.72553703362815e-08 wpclm = -2.9836416936794e-08 ppclm = 7.26033402456562e-15
+ pdiblc1 = 1.37328460825487 lpdiblc1 = -2.21762265468745e-07 wpdiblc1 = -1.28494787020665e-07 ppdiblc1 = 3.12676644840345e-14
+ pdiblc2 = 0.0418517851956429 lpdiblc2 = -7.49100245124536e-09 wpdiblc2 = -8.10624504834657e-09 ppdiblc2 = 1.97255745757456e-15
+ pdiblcb = 0.0440041723303621 lpdiblcb = -6.54589372865257e-08 wpdiblcb = -5.6982893580611e-07 ppdiblcb = 1.38661033581187e-13
+ drout = -0.975627884693997 ldrout = 3.42451386277089e-7
+ pscbe1 = 799752699.066856 lpscbe1 = 0.0428666491488912
+ pscbe2 = -6.28682802277113e-08 lpscbe2 = 1.7539304714853e-14 wpscbe2 = 6.3737152880367e-14 ppscbe2 = -1.55096713076027e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.97931790606873 lbeta0 = 5.63046413133249e-07 wbeta0 = 3.16208485163153e-06 pbeta0 = -7.69455403626315e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.86620788894034e-08 lagidl = -9.38361915278965e-15 wagidl = -3.43103089076314e-14 pagidl = 8.3490019489652e-21
+ bgidl = 1931628452.65062 lbgidl = -159.209155412696 wbgidl = 22.4408345339434 pbgidl = -5.46070779382105e-6
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0678392589988217 lkt1 = -1.08098220053745e-07 wkt1 = -1.1762176426676e-07 pkt1 = 2.86218448731447e-14
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080507e-08 wkt2 = -2.64697796016969e-23
+ at = 392704.922449648 lat = -0.0793644264910523 wat = -0.273858115484662 pat = 6.66400861058066e-8
+ ute = 0.608999778686825 lute = -1.93276019406095e-07 wute = -6.38637550815321e-07 pute = 1.55404784340299e-13
+ ua1 = 1.15501047585414e-09 lua1 = -1.83104660653394e-16 wua1 = -1.14202526933424e-16 pua1 = 2.77898144989255e-23
+ ub1 = -1.27707448617462e-19 lub1 = 1.37901457131676e-25 wub1 = 5.04223532089289e-25 pub1 = -1.22696745851543e-31
+ uc1 = 1.99309798377342e-10 luc1 = -4.83603756466256e-17 wuc1 = -1.77638117517771e-16 puc1 = 4.32261042405393e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.89 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.18282950331546 lvth0 = -1.52767356392756e-07 wvth0 = -4.81927361235598e-07 pvth0 = 8.6627619423399e-14
+ k1 = 2.87836403960321 lk1 = -2.15835788012492e-07 wk1 = -2.4585434495837e-06 pk1 = 3.48345952476648e-13
+ k2 = 0.332552009490551 lk2 = -9.93333847641458e-08 wk2 = -8.51286887496057e-08 pk2 = 1.98944414406093e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -115654.30229193 lvsat = -0.00430554846683723 wvsat = 0.273694675167753 pvsat = -1.62617383445883e-8
+ ua = -1.13210934489676e-08 lua = 1.17505946396009e-15 wua = 1.06916540095196e-14 pua = -1.49484028463845e-21
+ ub = -2.41049583718624e-18 lub = 7.34679397357211e-25 wub = 1.48312809221368e-24 pub = -1.97489777895946e-31
+ uc = 3.47186449884522e-12 luc = -4.70156804581691e-19 wuc = -2.56751950905138e-18 puc = 3.63254106313515e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0497138271649233 lu0 = 7.33915544591486e-09 wu0 = 5.26251830499949e-08 pu0 = -7.44632089008105e-15
+ a0 = -2.80402064513642 la0 = 5.46713443580799e-07 wa0 = 3.63093322898825e-06 pa0 = -5.15715656781089e-13
+ keta = -2.56245585355066 lketa = 4.28994291474924e-07 wketa = 2.0085560445651e-06 pketa = -3.30472705290292e-13
+ a1 = 0.0
+ a2 = -0.445070893740173 la2 = 2.07061902766929e-07 wa2 = -3.22323651831565e-07 pa2 = 4.62012276062329e-14
+ ags = 15.5143119325553 lags = -2.47254730176527e-06 wags = -9.83869789384694e-06 pags = 1.70542021552364e-12
+ b0 = 1.43374979148345e-05 lb0 = -2.48493431722792e-12 wb0 = -1.27566769372403e-11 pb0 = 2.21095092626587e-18
+ b1 = 1.61347698406525e-07 lb1 = -2.8012782434042e-14 wb1 = -1.43557856145158e-13 pb1 = 2.49241546709859e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -3.81298006685357 lvoff = 5.29312077260209e-07 wvoff = 2.83835366085893e-06 pvoff = -4.52578638091009e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -47.2436340978837 lnfactor = 7.30134576688018e-06 wnfactor = 3.90607490409127e-05 pnfactor = -5.38082319552591e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.170367210218553 leta0 = 5.95349459060933e-08 weta0 = -7.72138118459316e-07 peta0 = 8.71937434194953e-14
+ etab = 2.04177785855811 letab = -3.19135830065659e-07 wetab = -1.80239839608268e-06 petab = 2.76610674960542e-13
+ dsub = 0.560954466898676 ldsub = -4.55091431096207e-08 wdsub = -2.18998851535904e-07 pdsub = 3.35003753978878e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.12056326969416 lpclm = -8.87570992562366e-08 wpclm = 9.87921727200869e-07 ppclm = -1.69155827163968e-13
+ pdiblc1 = 0.28884401393627 lpdiblc1 = -3.37875017307465e-08 wpdiblc1 = 4.42765091483021e-07 ppdiblc1 = -6.77533803360373e-14
+ pdiblc2 = -0.013480476217546 lpdiblc2 = 2.10018107759398e-09 wpdiblc2 = 2.2066668515901e-08 ppdiblc2 = -3.25755503382498e-15
+ pdiblcb = -2.02861020764183 lpdiblcb = 2.93803894109094e-07 wpdiblcb = 1.41947856275986e-06 ppdiblcb = -2.06161549605241e-13
+ drout = 1.0
+ pscbe1 = 1457401859.61655 lpscbe1 = -113.952723542214 wpscbe1 = -453.330007749055 ppscbe1 = 7.85793168832055e-5
+ pscbe2 = 1.83190157256176e-07 lpscbe2 = -2.5111972721729e-14 wpscbe2 = -1.52143942285583e-13 ppscbe2 = 2.19107259662728e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 31.8017729021218 lbeta0 = -3.73962829097259e-06 wbeta0 = -1.39614869015835e-05 pbeta0 = 2.19871027693247e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.57054687871976e-08 lagidl = 8.70724282637701e-15 wagidl = 5.80339228614216e-14 pagidl = -7.65776249741889e-21
+ bgidl = 1075915243.7619 lbgidl = -10.8815392103429 wbgidl = -52.3619472458668 pbgidl = 7.50545679432816e-6
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.604058755002754 lkt1 = -1.51510050554153e-08 wkt1 = 2.74450783289105e-07 pkt1 = -3.93392263750941e-14
+ kt2 = -0.12
+ at = -136292.704278069 lat = 0.0123309641306765 wat = 0.335579971524386 pat = -3.89986930201676e-8
+ ute = -1.40013053483571 lute = 1.54982610879275e-07 wute = 1.03757183754526e-06 pute = -1.35145998619348e-13
+ ua1 = 1.16054941680031e-09 lua1 = -1.84064769599121e-16 wua1 = -7.16395182317985e-16 pua1 = 1.32172684997975e-22
+ ub1 = 2.09620272744075e-18 lub1 = -2.47586684965903e-25 wub1 = -1.17652157487501e-24 pub1 = 1.68640249499435e-31
+ uc1 = -4.98450921116467e-10 luc1 = 7.25880719489922e-17 wuc1 = 4.144889408748e-16 puc1 = -5.9412015807112e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.90 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0168761
+ k1 = 0.47866595
+ k2 = -0.0041430645
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 24491.02
+ ua = -9.0913219e-10
+ ub = 1.39839665e-18
+ uc = -6.8009552e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0102961633
+ a0 = 1.2509318
+ keta = 0.0074076058
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.23496304
+ b0 = -2.1309e-8
+ b1 = 2.2477e-9
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.34840646
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.0716757
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 790097310.0
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1731672e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.52561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.91 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.0168761
+ k1 = 0.47866595
+ k2 = -0.0041430645
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 24491.02
+ ua = -9.0913219e-10
+ ub = 1.39839665e-18
+ uc = -6.8009552e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0102961633
+ a0 = 1.2509318
+ keta = 0.0074076058
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.23496304
+ b0 = -2.1309e-8
+ b1 = 2.2477e-9
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.34840646
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.0716757
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 790097310.0
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1731672e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.52561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.92 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.08925744775245 lvth0 = 5.78568577480867e-7
+ k1 = 0.494917388074975 lk1 = -1.29903237519343e-7
+ k2 = -0.0325572332526668 lk2 = 2.27124054829104e-07 pk2 = 5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 13069.09495219 lvsat = 0.0912993075178117
+ ua = -9.66291472397079e-10 lua = 4.56893464037314e-16
+ ub = 2.21949209410947e-18 lub = -6.56329341502712e-24
+ uc = -6.33446214035016e-11 luc = -3.72883670043541e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0142698174381638 lu0 = -3.17627606214424e-8
+ a0 = 1.2538974524657 la0 = -2.37054625488884e-8
+ keta = 0.00418131295504559 lketa = 2.57888491967021e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.235883554325725 lags = -7.35798213936272e-9
+ b0 = -1.351101479895e-07 lb0 = 9.09651040668094e-13 wb0 = -2.52435489670724e-29
+ b1 = 4.795080260235e-09 lb1 = -2.03620714345863e-14 pb1 = -1.20370621524202e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.444837635940725 lvoff = 7.70806983031682e-07 wvoff = -4.2351647362715e-22
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 2.46027311128664 lnfactor = -3.10619045433921e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.395686193228354 lpclm = 3.17676376616597e-06 wpclm = 3.30872245021211e-24 ppclm = 3.91275008989622e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00124507074413753 lpdiblc2 = -3.2548529752527e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 780211112.930193 lpscbe1 = 79.0237147135631
+ pscbe2 = 9.45640285822898e-09 lpscbe2 = 4.90915183828849e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.78586633607361e-10 lalpha0 = -6.28169524705797e-16
+ alpha1 = 1.99833416432488e-10 lalpha1 = -7.98002241239631e-16
+ beta0 = -17.6314320251595 lbeta0 = 0.000164914009601124 wbeta0 = -6.7762635780344e-21
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.2445470400284e-09 lagidl = -8.56390118773294e-15
+ bgidl = 678903777.929449 lbgidl = 2566.63063353298
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.658049054769999 lkt1 = 1.05863012917712e-6
+ kt2 = -0.046450399725723 lkt2 = -4.82286063491885e-8
+ at = -42713.0729128486 lat = 0.421353408811043 pat = 1.05879118406788e-22
+ ute = -2.153658294925 lute = 7.14730947683921e-6
+ ua1 = -8.85759469220001e-10 lua1 = 5.03348062927607e-15
+ ub1 = 5.65236484917219e-19 lub1 = -5.6669956695524e-25
+ uc1 = 6.07016774048686e-11 luc1 = -4.19702820420277e-16 wuc1 = -1.23259516440783e-32 puc1 = 1.41059322098675e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.93 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.871079958408998 lvth0 = -2.92687881458923e-7
+ k1 = 0.475299486095559 lk1 = -5.15623240646724e-8
+ k2 = 0.040644405681078 lk2 = -6.51948315872987e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 39559.583135983 lvsat = -0.0144861655850803
+ ua = -1.08251348411575e-09 lua = 9.21007239869922e-16
+ ub = -8.03800002780308e-20 lub = 2.62087321463009e-24
+ uc = -7.89241966365168e-11 luc = 2.4926142797506e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00125238287902001 lu0 = 2.02202554661001e-8
+ a0 = 1.3338353970428 la0 = -3.42924694270506e-7
+ keta = 0.0265304661513564 lketa = -6.34588735299472e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.101537512133451 lags = 1.34007838455259e-6
+ b0 = 2.0447836173e-07 lb0 = -4.46440659558155e-13 pb0 = -1.92592994438724e-34
+ b1 = -9.64701613619999e-10 lb1 = 2.63868439399006e-15 wb1 = -3.94430452610506e-31
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.1977606647864 lvoff = -2.15854874803786e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.14967055274 lnfactor = 2.12748854560234e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.1392684955 letab = 2.76612515282979e-7
+ dsub = 0.859000699999999 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.498660454442519 lpclm = -3.94664687150745e-07 wpclm = 4.2351647362715e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00057063114206935 lpdiblc2 = -5.61587683608933e-10
+ pdiblcb = -0.424333799999999 lpdiblcb = 7.960072382244e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.63030196631712e-09 lpscbe2 = -2.03522732665583e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.87910516027147e-11 lalpha0 = -6.99185148545254e-17 walpha0 = -2.46519032881566e-32 palpha0 = 4.70197740328915e-38
+ alpha1 = 5.73670036880007e-16 lalpha1 = -2.15658830957128e-21 walpha1 = 9.4039548065783e-38 palpha1 = -6.27781712017518e-43
+ beta0 = 44.262864050319 lbeta0 = -8.22508349003348e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.5111712326491e-10 lagidl = 1.00279555078445e-15
+ bgidl = 1642192444.1411 lbgidl = -1280.10660221933
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.29548101427894 lkt1 = -3.89226604501367e-7
+ kt2 = -0.0595514414067929 lkt2 = 4.08828123541189e-9
+ at = 85592.4759078148 lat = -0.0910140149053682
+ ute = 0.23572003740572 lute = -2.39428581403369e-6
+ ua1 = 7.57014667690222e-10 lua1 = -1.52667175706473e-15
+ ub1 = 3.3072320827312e-19 lub1 = 3.69791212172155e-25
+ uc1 = -1.34630329173249e-10 luc1 = 3.6032390406437e-16 wuc1 = 4.93038065763132e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.94 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.049504128414 lvth0 = 6.29717967305065e-8
+ k1 = 0.414136178847399 lk1 = 7.03568204787615e-8
+ k2 = 0.019004695517398 lk2 = -2.20595750090491e-08 wk2 = -1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -120709.932052356 lvsat = 0.304985149281413 pvsat = 5.29395592033938e-23
+ ua = -2.38835009088599e-10 lua = -7.60729124183748e-16
+ ub = 1.22011089563328e-18 lub = 2.85552931560295e-26
+ uc = -1.0751845924825e-10 luc = 8.1924173043452e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0140859613026 lu0 = -5.3614040816021e-09 wu0 = -1.32348898008484e-23
+ a0 = 1.1025970552 la0 = 1.18011479581738e-7
+ keta = -0.0111645336712126 lketa = 1.16800020263728e-8
+ a1 = 0.0
+ a2 = 1.1973352 la2 = -7.920233528976e-7
+ ags = 0.68894229203862 lags = -2.35615047336159e-7
+ b0 = -1.61612814364e-07 lb0 = 2.83302793214707e-13 pb0 = -7.22223729145213e-35
+ b1 = 2.8206905647e-09 lb1 = -4.90688167995797e-15 wb1 = 7.88860905221012e-31 pb1 = 3.76158192263132e-37
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.35231008046714 lvoff = 9.22143483504274e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -0.341843953883803 lnfactor = 5.10058108920683e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.485738951 leta0 = 9.69238578108438e-07 weta0 = -1.57164316385075e-22 peta0 = -2.20881053461883e-29
+ etab = 0.162904101 letab = -3.25719603879139e-07 wetab = 5.12851979782877e-23 petab = 2.20881053461883e-29
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0742494148848616 lpclm = 7.47338325954558e-7
+ pdiblc1 = 0.389494937293899 lpdiblc1 = 1.00676068445305e-9
+ pdiblc2 = 0.000148737715861299 lpdiblc2 = 2.79388514801769e-10
+ pdiblcb = 0.1736676 lpdiblcb = -3.960116764488e-07 ppdiblcb = -1.51461293802434e-28
+ drout = 0.233817461872679 ldrout = 6.50192048185637e-7
+ pscbe1 = 801195690.883978 lpscbe1 = -2.38341607528855
+ pscbe2 = 1.00453763670072e-08 lpscbe2 = -1.03090630838839e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.19286376348734e-11 lalpha0 = 1.9065000905095e-16 walpha0 = -6.16297582203915e-33 palpha0 = -5.87747175411144e-39
+ alpha1 = -9.93348130700257e-11 lalpha1 = 1.98006844545353e-16 walpha1 = -5.91922531345265e-33 palpha1 = 8.26497941477509e-38
+ beta0 = -1.89174393923941 lbeta0 = 9.75089908035558e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.57762120486598e-11 lagidl = 5.50520443557167e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.46303225874108 lkt1 = -5.52403419676924e-8
+ kt2 = -0.0552956877620159 lkt2 = -4.39487422336052e-9
+ at = 7282.96884286986 lat = 0.0650833012884552
+ ute = -1.74526153944298 lute = 1.55448004039875e-6
+ ua1 = -1.01421246704804e-09 lua1 = 2.00398259724017e-15 wua1 = -7.39557098644699e-32 pua1 = -3.76158192263132e-37
+ ub1 = 1.51236168895956e-18 lub1 = -1.98561367364239e-24 wub1 = -7.3468396926393e-40
+ uc1 = 9.45390689071462e-11 luc1 = -9.64881655664091e-17 puc1 = 4.70197740328915e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.95 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.021185345124 lvth0 = 3.48416731747835e-8
+ k1 = 0.433942827763722 lk1 = 5.06821234575217e-8
+ k2 = 0.0053098971143308 lk2 = -8.45601135294313e-09 pk2 = -3.15544362088405e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 281821.671312781 lvsat = -0.0948647885421043
+ ua = -2.19856609529999e-10 lua = -7.79581089644489e-16
+ ub = 6.40974805810801e-19 lub = 6.03833178348113e-25
+ uc = -3.68425960659401e-11 luc = 1.17191524616627e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0119524255404 lu0 = -3.24208193464985e-9
+ a0 = 1.3370384272 la0 = -1.14868043997993e-7
+ keta = 0.0102543614029353 lketa = -9.59620036879108e-09 wketa = 1.65436122510606e-24 pketa = -1.57772181044202e-30
+ a1 = 0.0
+ a2 = 0.00532960000000049 la2 = 3.920411057952e-7
+ ags = 0.0750739951768802 lags = 3.74163658931889e-7
+ b0 = 2.21467272524e-07 lb0 = -9.72252141344452e-14
+ b1 = -2.05039325756e-08 lb1 = 1.82623528209814e-14 wb1 = 3.15544362088405e-30 pb1 = 3.00926553810506e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.17299845369812 lvoff = -8.59027043610566e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 7.20701764227201 lnfactor = -2.39798999099538e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -0.327795373275 letab = 1.61710830498242e-7
+ dsub = 0.22285388835452 ldsub = 3.68986442496979e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.724860464581081 lpclm = -4.64478834943812e-8
+ pdiblc1 = 0.582254436329561 lpdiblc1 = -1.90468574568633e-07 wpdiblc1 = 4.2351647362715e-22
+ pdiblc2 = -6.97233132010396e-05 lpdiblc2 = 4.96394156488494e-10
+ pdiblcb = -0.225
+ drout = 0.940647677979241 ldrout = -5.19292650212225e-8
+ pscbe1 = 797608618.23204 lpscbe1 = 1.17975949864194
+ pscbe2 = 1.69084195225236e-08 lpscbe2 = -7.84822787040275e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.80525548816681 lbeta0 = 1.11183906313476e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.2751125890816e-10 lagidl = -2.95540344420154e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.527763005202081 lkt1 = 9.05916826038275e-9
+ kt2 = -0.0440516586270121 lkt2 = -1.55639956362672e-8
+ at = 79613.5535857882 lat = -0.00676541709890555
+ ute = -0.267515207816925 lute = 8.65784548339858e-8
+ ua1 = 1.6847864446152e-09 lua1 = -6.77035583673575e-16
+ ub1 = -1.43727939498936e-18 lub1 = 9.44376901405261e-25 pub1 = -3.50324616081204e-46
+ uc1 = -2.91537921926444e-11 luc1 = 2.63806536927348e-17 wuc1 = 6.16297582203915e-33 puc1 = 1.0285575569695e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.96 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.939594243016002 lvth0 = -5.41031795697235e-9
+ k1 = 0.494267157497442 lk1 = 2.09218392753482e-8
+ k2 = -0.00919181642799757 lk2 = -1.30176499739792e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67329.9919879199 lvsat = 0.0109521075526635
+ ua = -2.0449807407592e-09 lua = 1.20821999007862e-16
+ ub = 2.041231234016e-18 lub = -8.69665274297851e-26
+ uc = -2.58807559379872e-11 luc = 6.31126017661872e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00522382485816002 lu0 = 7.73924687250611e-11
+ a0 = 1.38850638568 la0 = -1.402591436986e-7
+ keta = -0.008445362407908 lketa = -3.7091602339729e-10
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = 1.23423871552472 lags = -1.97696345875074e-7
+ b0 = 4.8132028632e-08 lb0 = -1.17123515832536e-14
+ b1 = 3.2587934928e-08 lb1 = -7.92988290950966e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.2740601181368 lvoff = -3.60451449502073e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 1.68816362963119 lnfactor = 3.24670409892803e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 4.850105e-05 letab = -2.70107735049e-11 petab = 3.08148791101958e-33
+ dsub = -0.023901594981119 ldsub = 1.58632500887536e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.624438894129922 lpclm = 3.09389322885369e-9
+ pdiblc1 = -0.0625215999738398 lpdiblc1 = 1.27623945629214e-07 ppdiblc1 = -5.04870979341448e-29
+ pdiblc2 = -0.0089245210323659 lpdiblc2 = 4.86480235366586e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = -7.88860905221012e-31
+ pdiblcb = -0.225
+ drout = 1.22833572426512 ldrout = -1.93856710399806e-07 wdrout = 8.470329472543e-22
+ pscbe1 = 800069244.26128 lpscbe1 = -0.0341608253716004
+ pscbe2 = -6.99090056320879e-09 lpscbe2 = 3.9422149020523e-15 ppscbe2 = -1.1284745767894e-36
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.83100208558321 lbeta0 = 1.12461288258562e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.5080962010832e-10 lagidl = -1.09699111337918e-16
+ bgidl = 730034204.006401 lbgidl = 133.18438586389
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.50680115016 lkt1 = -1.28211138236603e-9
+ kt2 = -0.132062202816 lkt2 = 2.78549502128398e-8
+ at = 65261.4810880001 lat = 0.000315005643008265
+ ute = -0.0012549260000001 lute = -4.47778600770119e-8
+ ua1 = 2.2472125128e-10 lua1 = 4.32700586760273e-17
+ ub1 = 5.1394790896e-19 lub1 = -1.82376742705086e-26
+ uc1 = 4.74348323563201e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.97 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.772463663771422 lvth0 = -4.60795388491882e-8
+ k1 = -0.41547953916943 lk1 = 2.4229778094887e-7
+ k2 = 0.438589349394086 lk2 = -1.10263938326212e-07 wk2 = 5.29395592033938e-23 pk2 = 4.41762106923767e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 92623.7868717136 lvsat = 0.00479716609323066
+ ua = -1.55915274021428e-09 lua = 2.60158501126276e-18
+ ub = 9.27892317999923e-20 lub = 3.87163452505452e-25
+ uc = 6.09622494694269e-15 luc = 1.20053449946549e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00281915098371424 lu0 = 6.62540999984932e-10
+ a0 = -0.397764477428577 la0 = 2.94408435588514e-7
+ keta = -0.184161871607297 lketa = 4.23875878921637e-08 wketa = 2.64697796016969e-23 pketa = -6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.164955374457998 la2 = 8.73018597320191e-8
+ ags = -1.62902379023886 lags = 4.99044225752424e-07 pags = 2.01948391736579e-28
+ b0 = 1.23812857142857e-09 lb0 = -3.01283730314285e-16
+ b1 = -1.86798933828571e-10 lb1 = 4.54552789599769e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.403685441391142 lvoff = -4.50237804014223e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -5.5978371627743 lnfactor = 2.09763127071517e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.39713389074943 leta0 = -2.20740146707184e-7
+ etab = 0.244655617911143 letab = -5.95492173762616e-08 wetab = 1.6130021944784e-23 petab = -1.1339875512552e-29
+ dsub = 1.53653693089571 ldsub = -2.21081489122281e-07 pdsub = 2.01948391736579e-28
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.664807054980852 lpclm = -6.72921429629145e-9
+ pdiblc1 = 1.18699067550629 lpdiblc1 = -1.76429872461569e-7
+ pdiblc2 = 0.0300992129326342 lpdiblc2 = -4.63115502190936e-09 wpdiblc2 = -2.64697796016969e-23
+ pdiblcb = -0.78214353300956 lpdiblcb = 1.35574193035481e-7
+ drout = -0.975627884694001 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066856 lpscbe1 = 0.0428666491488912
+ pscbe2 = 2.95389305828886e-08 lpscbe2 = -4.94688114937674e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 11.56376242988 lbeta0 = -5.52523148401942e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.10815918728486e-08 lagidl = 2.72090620315522e-15 wagidl = 2.76101316827354e-30 pagidl = 4.70197740328915e-37
+ bgidl = 1964163557.12 lbgidl = -167.126182664067
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.238369297999997 lkt1 = -6.66017814232763e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080508e-08 wkt2 = -5.29395592033938e-23 pkt2 = -2.52435489670724e-29
+ at = -4339.24200000009 lat = 0.017251506397796
+ ute = -0.316907829714285 lute = 3.20324862070149e-8
+ ua1 = 9.8943770542857e-10 lua1 = -1.42814513843578e-16 wua1 = 7.88860905221012e-31
+ ub1 = 6.03324423999999e-19 lub1 = -3.9986376687312e-26
+ uc1 = -5.82329727011429e-11 luc1 = 1.43095671820707e-17 wuc1 = -2.31111593326468e-32 puc1 = 3.67341984631965e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.98 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.520352091175162 lvth0 = -8.97800546198801e-08 wvth0 = -2.49123788935557e-07 pvth0 = 4.31826193265113e-14
+ k1 = -4.11333191723232 lk1 = 8.83276116457536e-07 wk1 = 2.36392430141515e-06 pk1 = -4.097579105587e-13
+ k2 = 1.33266162872819 lk2 = -2.65240639081427e-07 wk2 = -7.74946497763736e-07 pk2 = 1.3432767602937e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 553155.212815385 lvsat = -0.0750304302169931 wvsat = -0.187611471163299 pvsat = 3.25201971885039e-8
+ ua = 1.02679182791027e-08 lua = -2.04747925133511e-15 wua = -4.19919843562542e-15 pua = 7.27880658434437e-22
+ ub = -4.24535660405064e-18 lub = 1.13912897540013e-24 wub = 2.74870899424445e-24 pub = -4.76455719644343e-31
+ uc = 2.07223916932761e-13 luc = -2.2857726878783e-20 wuc = -3.15759131873796e-19 puc = 5.47330564007401e-26
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0444091931970076 lu0 = -6.5465937371829e-09 wu0 = -1.22954360850881e-08 pu0 = 2.13126630011701e-15
+ a0 = -10.6730705149987 la0 = 2.07550943352884e-06 wa0 = 9.05854899813677e-06 pa0 = -1.57019076623903e-12
+ keta = -0.441264945469912 lketa = 8.69533205093617e-08 wketa = 5.45481161005485e-07 pketa = -9.45526134863688e-14
+ a1 = 0.0
+ a2 = -7.2643021704831 la2 = 1.37507450405702e-06 wa2 = 4.38118793129792e-06 pa2 = -7.59426353635319e-13
+ ags = 21.1495017276852 lags = -3.4493398304735e-06 wags = -1.37255261005574e-05 pags = 2.37915524321842e-12
+ b0 = -1.01826005104488e-05 lb0 = 1.76494493828017e-12 wb0 = 4.15586969483117e-12 pb0 = -7.20370141162646e-19
+ b1 = 3.81162611686897e-07 lb1 = -6.60568888592154e-14 wb1 = -2.95173478023971e-13 pb1 = 5.11647803337191e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 4.55595098084441 lvoff = -8.64195836197608e-07 wvoff = -2.93405125162859e-06 pvoff = 5.08582575854796e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 8.69002721260188 lnfactor = -3.78998564383784e-07 wnfactor = 4.80942434563544e-07 pnfactor = -8.33655997223732e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -6.31559897469831 leta0 = 1.1161695427238e-06 weta0 = 3.70150646705085e-06 peta0 = -6.4161172798566e-13
+ etab = -1.28158713182753 letab = 2.05006648377941e-07 wetab = 4.89866683788896e-07 petab = -8.49125112345996e-14
+ dsub = 0.0907377406737719 ldsub = 2.95304509124099e-08 wdsub = 1.0532946768726e-07 pdsub = -1.82575992699743e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 15.1235848598275 lpclm = -2.5129848414328e-06 wpclm = -8.6705531910252e-06 ppclm = 1.50293634902593e-12
+ pdiblc1 = 6.28425096755649 lpdiblc1 = -1.05997877696497e-06 wpdiblc1 = -3.69252009060229e-06 ppdiblc1 = 6.4005404746482e-13
+ pdiblc2 = 0.127385736727115 lpdiblc2 = -2.1494606483397e-08 wpdiblc2 = -7.5094703106218e-08 ppdiblc2 = 1.30167656470256e-14
+ pdiblcb = -2.16260086989224 lpdiblcb = 3.7485990689605e-07 wpdiblcb = 1.51189757691991e-06 ppdiblcb = -2.62069302188144e-13
+ drout = 1.0
+ pscbe1 = 801197746.521767 lpscbe1 = -0.207614986587942 wpscbe1 = -0.718339133996778 ppscbe1 = 1.24515468808914e-7
+ pscbe2 = -2.57115376447668e-08 lpscbe2 = 4.6301245122686e-15 wpscbe2 = -8.0556276608785e-15 ppscbe2 = 1.39634638748135e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.1646409435277 lbeta0 = -8.30016228200577e-07 wbeta0 = -1.10667050277243e-06 pbeta0 = 1.91828051609566e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.17461625048231e-08 lagidl = -1.23601108516162e-15 wagidl = 4.61226430047438e-15 pagidl = -7.99480669315629e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 1.93948854361926 lkt1 = -4.44107303973876e-07 wkt1 = -1.4799411262665e-06 pkt1 = 2.56530034944782e-13
+ kt2 = -0.12
+ at = 886727.42584506 lat = -0.137204207673131 wat = -0.370040183671028 pat = 6.41420253571686e-8
+ ute = 5.88488445721897 lute = -1.04297378522542e-06 wute = -3.98721043010752e-06 pute = 6.91135081533978e-13
+ ua1 = -6.25358620211367e-10 lua1 = 1.37091051650198e-16 wua1 = 5.15420956128132e-16 pua1 = -8.9342037693338e-23
+ ub1 = 5.09221917644162e-19 lub1 = -2.36748364406034e-26 wub1 = -8.19139397681272e-26 pub1 = 1.41987984915277e-32
+ uc1 = 6.3301884706147e-10 luc1 = -1.05510640751941e-16 wuc1 = -3.65933506261741e-16 puc1 = 6.34301821083976e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.99 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.13181153747554 wvth0 = 6.89316321295417e-8
+ k1 = 0.5536725055272 wk1 = -4.49845966263051e-8
+ k2 = -0.0764006435052808 wk2 = 4.33359193993009e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -248939.518899277 wvsat = 0.163987832946638
+ ua = -1.34314287141275e-09 wua = 2.60294520893984e-16
+ ub = 4.39741842647386e-18 wub = -1.79863991807034e-24
+ uc = -4.87091391354924e-12 wuc = -3.78669057109717e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.022432676439988 wu0 = -7.27877909090531e-9
+ a0 = 0.0081446176441542 wa0 = 7.45351918877897e-7
+ keta = -0.0550604796320326 wketa = 3.74647469867952e-8
+ a1 = 0.0
+ a2 = 0.0791263930769226 wa2 = 4.32338322937981e-7
+ ags = 0.592480648626646 wags = -2.14418397136484e-7
+ b0 = -6.29827212832308e-08 wb0 = 2.49934892845916e-14
+ b1 = 1.41734032646154e-09 wb1 = 4.98001737399239e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.425953345210784 wvoff = 4.65081395394634e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 3.15617132384077 wnfactor = -6.50417791332635e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.00752026452741314 wpclm = -3.46652798468104e-9
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00486236335036257 wpdiblc2 = 3.41867350676308e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1313834677.59128 wpscbe1 = -314.107401061401
+ pscbe2 = 8.13931185585953e-09 wpscbe2 = 8.26748547497198e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.61340153846154e-10 walpha0 = -2.16710938816031e-16
+ alpha1 = 4.61340153846154e-10 walpha1 = -2.16710938816031e-16
+ beta0 = -94.5618415384615 wbeta0 = 5.85119534803283e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.37464993751129e-09 wagidl = -1.32032210025704e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.20164129383077 wkt1 = 4.05444495430912e-7
+ kt2 = -0.0291177113072416 wkt2 = -1.40137493864301e-8
+ at = -261141.0696175 wat = 0.162614741602753
+ ute = -4.72388485901538 wute = 2.07773779699258e-6
+ ua1 = -3.41965361665512e-09 wua1 = 1.8973465929807e-15
+ ub1 = 1.39510181602126e-18 wub1 = -5.40224873216586e-25
+ uc1 = -2.12165063617345e-10 wuc1 = 1.32159289320226e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.100 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.097385963809 lvth0 = -6.8828213015911e-07 wvth0 = 4.82851628425066e-08 pvth0 = 4.12791838962311e-13
+ k1 = 0.578425765536448 lk1 = -4.94900293966763e-07 wk1 = -5.98301712414229e-08 pk1 = 2.96812591084273e-13
+ k2 = -0.062650490227771 lk2 = -2.7491146202906e-07 wk2 = 3.508937222231e-08 pk2 = 1.64876005042525e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -390400.785728908 lvsat = 2.82828292163301 wvsat = 0.248828124329828 pvsat = -1.69624062164261e-6
+ ua = -1.34647393985968e-09 lua = 6.6599177360481e-17 wua = 2.62292303212693e-16 pua = -3.9942337148363e-23
+ ub = 4.36537977955187e-18 lub = 6.40559496973946e-25 wub = -1.77942498948033e-24 pub = -3.84170561946047e-31
+ uc = 6.18083202565629e-12 luc = -2.20961292052666e-16 wuc = -4.4495104134392e-17 puc = 1.32519811410508e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0225016375839453 lu0 = -1.37876346000426e-09 wu0 = -7.32013799909675e-09 pu0 = 8.26902630782492e-16
+ a0 = -0.780226219859202 la0 = 1.57621646235477e-05 wa0 = 1.218171179378e-06 pa0 = -9.45323528808866e-12
+ keta = -0.0903377472911431 lketa = 7.05310336025064e-07 wketa = 5.8622013102659e-08 pketa = -4.23004372610411e-13
+ a1 = 0.0
+ a2 = -0.401055806541017 la2 = 9.60044501854497e-06 wa2 = 7.20323851737685e-07 pa2 = -5.7577920164012e-12
+ ags = 0.80716748652396 lags = -4.29230651423221e-06 wags = -3.43175153608062e-07 pags = 2.57427735191996e-12
+ b0 = 3.03751078259463e-07 lb0 = -7.33223281028131e-12 wb0 = -1.94952246467502e-13 pb0 = 4.3974494365503e-18
+ b1 = -1.17892346664391e-08 lb1 = 2.6404351765541e-13 wb1 = 8.41854207810647e-15 pb1 = -1.58358040174395e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.284051562360231 lvoff = -2.83709030733373e-06 wvoff = -3.85963478912499e-08 pvoff = 1.70152278251901e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 3.40491942273428 lnfactor = -4.97330481803539e-06 wnfactor = -7.99602523408848e-07 pnfactor = 2.98270077283915e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.03464159443462e-06 lcit = 2.4061265710639e-10 wcit = 7.21768242605774e-12 pcit = -1.44305564320832e-16
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.48248108775496 lpclm = -2.94893902755465e-05 wpclm = -8.88062777020979e-07 ppclm = 1.76860318005149e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00947587760059476 lpdiblc2 = 9.22395497727087e-08 wpdiblc2 = 6.18559269292869e-09 ppdiblc2 = -5.53199505076938e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1656546466.01729 lpscbe1 = -6851.95262258565 wpscbe1 = -519.646123017949 ppscbe1 = 0.00410940514016528
+ pscbe2 = 7.14432644037761e-09 lpscbe2 = 1.98930797168004e-14 wpscbe2 = 1.42348328954624e-15 ppscbe2 = -1.19307193941293e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.02032985734846e-10 lalpha0 = -4.8122531421278e-15 walpha0 = -3.61064587337185e-16 palpha0 = 2.88611128641664e-21
+ alpha1 = 7.02032985734846e-10 lalpha1 = -4.8122531421278e-15 walpha1 = -3.61064587337185e-16 palpha1 = 2.88611128641664e-21
+ beta0 = -155.154652694166 lbeta0 = 0.00121145255380617 wbeta0 = 9.4852019347035e-05 pbeta0 = -7.26559219815329e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.04976259448444e-09 lagidl = -1.34977555389422e-14 wagidl = -1.72521565039797e-15 pagidl = 8.0951736019874e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.32198770977512 lkt1 = 2.4061265710639e-06 wkt1 = 4.77621319691489e-07 pkt1 = -1.44305564320832e-12
+ kt2 = -0.0291177113072416 wkt2 = -1.40137493864301e-8
+ at = -261141.0696175 wat = 0.162614741602753
+ ute = -4.72388485901539 wute = 2.07773779699258e-6
+ ua1 = -3.41965361665512e-09 wua1 = 1.8973465929807e-15
+ ub1 = 1.39510181602126e-18 wub1 = -5.40224873216587e-25
+ uc1 = -2.28532176185776e-10 luc1 = 3.2723321366469e-16 wuc1 = 1.41975337419665e-16 puc1 = -1.96255567476332e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.101 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.75153208386546 lvth0 = 4.5405289088408e-06 wvth0 = 3.97194047266617e-07 pvth0 = -2.37615480544253e-12
+ k1 = 0.591486079244702 lk1 = -5.99295795822876e-07 wk1 = -5.79163192932525e-08 pk1 = 2.81514525580591e-13
+ k2 = -0.306675478305555 lk2 = 1.67566274812264e-06 wk2 = 1.64400279348158e-07 pk2 = -8.68749782700989e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -89264.695165759 lvsat = 0.421200365763145 wvsat = 0.061373892419677 pvsat = -1.97855586454384e-7
+ ua = -1.56280940607658e-09 lua = 1.79584168021972e-15 wua = 3.57756977884394e-16 pua = -8.03023748859311e-22
+ ub = 1.05062939588489e-17 lub = -4.84458431671395e-23 wub = -4.9699447813229e-24 pub = 2.51187325299413e-29
+ uc = 5.88486504932358e-14 luc = -1.72026209704606e-16 wuc = -3.80257366178169e-17 puc = 8.08079702043027e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.052594110308384 lu0 = -2.41918069202224e-07 wu0 = -2.29846957194301e-08 pu0 = 1.26039007109917e-13
+ a0 = 1.20536821402319 la0 = -1.09362817392919e-07 wa0 = 2.91050322278374e-08 pa0 = 5.13723304403464e-14
+ keta = -0.0169846600745327 lketa = 1.18974316559218e-07 wketa = 1.26941272299e-08 pketa = -5.58872572040236e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.274428699785491 lags = -3.3945326121706e-08 wags = -2.31171503373601e-08 pags = 1.59455521721278e-14
+ b0 = -1.836440293434e-06 lb0 = 9.77504020834815e-12 wb0 = 1.0203594843552e-12 pb0 = -5.31694800328061e-18
+ b1 = 4.80223568679698e-08 lb1 = -2.14050749797058e-13 wb1 = -2.59252219727314e-14 pb1 = 1.16163274076201e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -1.35203925379799 lvoff = 5.69969629016802e-06 wvoff = 5.44087094137278e-07 pvoff = -2.95606291661842e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 6.14613801227154 lnfactor = -2.688479153609e-05 wnfactor = -2.21056872461946e-06 pnfactor = 1.42610305256916e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.80670076923077e-05 wcit = -1.08355469408015e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.04025260894415 lpclm = 1.46556868461589e-05 wpclm = 2.18580028020751e-06 ppclm = -6.88439458162576e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00394223301804862 lpdiblc2 = -1.50159437234969e-08 wpdiblc2 = -1.61760203591244e-09 ppdiblc2 = 7.05362243975163e-15
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 753729551.529228 lpscbe1 = 364.56812703449 wpscbe1 = 15.8821098940512 ppscbe1 = -0.00017125303404306
+ pscbe2 = 9.34969932120297e-09 lpscbe2 = 2.26478886432963e-15 wpscbe2 = 6.39946140437645e-17 ppscbe2 = -1.06386690366568e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.62551696386713e-10 lalpha0 = -2.89799825169237e-15 walpha0 = -1.70305831474426e-16 palpha0 = 1.36131207434613e-21
+ alpha1 = 5.60571636959512e-10 lalpha1 = -3.68150476743067e-15 walpha1 = -2.16349934002962e-16 palpha1 = 1.72935814876337e-21
+ beta0 = -98.7779539734964 lbeta0 = 0.000760814545607688 wbeta0 = 4.86669935956439e-05 pbeta0 = -3.57386698445756e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.30384235137417e-09 lagidl = -3.95087149147197e-14 wagidl = -3.0342729004762e-15 pagidl = 1.85589106632132e-20
+ bgidl = -481345804.894464 lbgidl = 11840.8977134035 wbgidl = 695.850637351896 pbgidl = -0.00556216934186913
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.69426959642841 lkt1 = 5.38190152236133e-06 wkt1 = 6.21465187339403e-07 pkt1 = -2.59284829654537e-12
+ kt2 = 0.011922586986256 lkt2 = -3.28048975880749e-07 wkt2 = -3.50087434712131e-08 pkt2 = 1.67820084027671e-13
+ at = -580986.793542041 lat = 2.55663497918354 wat = 0.322825465412337 pat = -1.28061846663466e-6
+ ute = -10.1128068191824 lute = 4.30754746832378e-05 wute = 4.77343724606491e-06 pute = -2.1547636842849e-11
+ ua1 = -8.66252479772217e-09 lua1 = 4.19080414407281e-14 wua1 = 4.66405434699961e-15 pua1 = -2.2115230225094e-20
+ ub1 = 3.43513366812909e-18 lub1 = -1.63066641246639e-23 wub1 = -1.72119845043329e-24 pub1 = 9.43992097176223e-30
+ uc1 = -1.23024314965974e-11 luc1 = -1.40116422128962e-15 wuc1 = 4.37836448816047e-17 puc1 = 5.8862381977246e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.102 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.244253887818843 lvth0 = -1.47854238800361e-06 wvth0 = -3.75934046593098e-07 pvth0 = 7.1120699063503e-13
+ k1 = 0.420797466108852 lk1 = 8.23215291798104e-08 wk1 = 3.26871613712719e-08 pk1 = -8.02957966893227e-14
+ k2 = 0.221708244813498 lk2 = -4.34352051990156e-07 wk2 = -1.08591625221724e-07 pk2 = 2.21399163510295e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 61722.9094512185 lvsat = -0.181744173282808 wvsat = -0.0132922820836173 pvsat = 1.00311685504252e-7
+ ua = -2.01297051172557e-09 lua = 3.59348712952987e-15 wua = 5.58034344744174e-16 pua = -1.60279896848041e-21
+ ub = -4.21144103905679e-18 lub = 1.03270472739271e-23 wub = 2.47757163573146e-24 pub = -4.62171778390572e-30
+ uc = -5.38300131134682e-11 luc = 4.31702297541683e-17 wuc = -1.5050040833317e-17 puc = -1.09417488483803e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0273162283959642 lu0 = 7.71909229387209e-08 wu0 = 1.71338017770039e-08 pu0 = -3.41677134454981e-14
+ a0 = 1.54668355629703 la0 = -1.47235034367806e-06 wa0 = -1.27654023297083e-07 pa0 = 6.77364223712119e-13
+ keta = 0.0581517503400803 lketa = -1.81070766333052e-07 wketa = -1.89646185461705e-08 pketa = 7.05368153358982e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.769227313045396 lags = 4.13372588884437e-06 wags = 4.00441750116493e-07 pags = -1.67546830024846e-12
+ b0 = 1.22393762790181e-06 lb0 = -2.44608323928315e-12 wb0 = -6.11412743104268e-13 pb0 = 1.19927003997794e-18
+ b1 = 1.16548799309345e-08 lb1 = -6.88231221802718e-14 wb1 = -7.56849559861051e-15 pb1 = 4.28586610908223e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.315997186170879 lvoff = -9.61337010944397e-07 wvoff = -3.0812226380039e-07 pvoff = 4.4709709638967e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -3.10848396148035 lnfactor = 1.00720420673285e-05 wnfactor = 2.55379495629844e-06 pnfactor = -4.76468400713777e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.80670076923077e-05 wcit = -1.08355469408015e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.1592351855 leta0 = -3.16412877194199e-7
+ etab = -0.1392684955 letab = 2.76612515282979e-7
+ dsub = 0.8590007 ldsub = -1.1940108573366e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0251475491022051 lpclm = -1.57883009017358e-06 wpclm = 2.83985671577193e-07 ppclm = 7.10193963972804e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00362348161614442 lpdiblc2 = -1.37430616377196e-08 wpdiblc2 = -1.83092325959283e-09 ppdiblc2 = 7.90548618848105e-15
+ pdiblcb = -1.14460685958738 lpdiblcb = 3.67230101745096e-06 wpdiblcb = 4.31978149357668e-07 ppdiblcb = -1.72503475899965e-12
+ drout = 0.56
+ pscbe1 = 889897293.439555 lpscbe1 = -179.195691110215 wpscbe1 = -53.9152005414844 ppscbe1 = 0.000107471218016962
+ pscbe2 = 1.00279120245314e-08 lpscbe2 = -4.43543695954518e-16 wpscbe2 = -2.3846353105557e-16 ppscbe2 = 1.43950700569001e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.4251798649734e-10 lalpha0 = 1.11558470561647e-15 walpha0 = 3.48635561390011e-16 palpha0 = -7.10996309552359e-22
+ alpha1 = -7.21474037069614e-10 lalpha1 = 1.43813694040546e-15 walpha1 = 4.32698770289142e-16 palpha1 = -8.62512705937055e-22
+ beta0 = 277.427250265833 lbeta0 = -0.00074149999227899 wbeta0 = -0.000139838521950542 pbeta0 = 3.95379539994421e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.23641794250093e-09 lagidl = 6.57544504670294e-15 wagidl = 2.45012730099042e-15 pagidl = -3.34215306851105e-21
+ bgidl = 3962691609.78892 lbgidl = -5905.64576807343 wbgidl = -1391.70127470379 pbgidl = 0.0027741310355155
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.07695428438333 lkt1 = -1.07658517121012e-06 wkt1 = -1.31059701746399e-07 pkt1 = 4.12237938986756e-13
+ kt2 = -0.0749495632854872 lkt2 = 1.8860882941113e-08 wkt2 = 9.23490349139609e-09 pkt2 = -8.85975264670087e-15
+ at = 201781.238246617 lat = -0.569222347343314 wat = -0.0696833039403501 pat = 2.86801717354665e-7
+ ute = 2.85389809823818 lute = -8.70496079828483e-06 wute = -1.5702318701954e-06 pute = 3.78477809853975e-12
+ ua1 = 3.59568907585836e-09 lua1 = -7.04314983276821e-15 wua1 = -1.70247283463846e-15 pua1 = 3.30846469737417e-21
+ ub1 = -1.07554373303467e-18 lub1 = 1.70599534714458e-24 wub1 = 8.43397629167203e-25 pub1 = -8.01378007557458e-31
+ uc1 = -7.79450885908582e-10 luc1 = 1.66231885335503e-15 wuc1 = 3.86726099301673e-16 puc1 = -7.80861315276469e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.103 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -1.05323975815205 lvth0 = 1.34039888794637e-07 wvth0 = 2.24041479748154e-09 pvth0 = -4.26225338843454e-14
+ k1 = 0.296664741042692 lk1 = 3.2976000709774e-07 wk1 = 7.04525785461585e-08 pk1 = -1.55575037829876e-13
+ k2 = 0.0594185680367042 lk2 = -1.10853872263255e-07 wk2 = -2.42379048152482e-08 pk2 = 5.32536871826916e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -736385.081480147 lvsat = 1.40915481314434 wvsat = 0.369246368603152 pvsat = -6.62217143378412e-7
+ ua = -1.11166001428523e-10 lua = -1.97452069416628e-16 wua = -7.65684915258714e-17 pua = -3.37821020035555e-22
+ ub = 1.62103739275318e-18 lub = -1.29905361838012e-24 wub = -2.40452539420981e-25 pub = 7.96223089344296e-31
+ uc = -1.09088769677893e-10 luc = 1.53319609046787e-16 wuc = 9.41781431757296e-19 puc = -4.28188558585991e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0142690965237155 lu0 = -5.70268546602359e-09 wu0 = -1.09833920409283e-10 pu0 = 2.04680848312011e-16
+ a0 = -0.657346400237806 la0 = 2.92102632182118e-06 wa0 = 1.05551235983987e-06 pa0 = -1.68108628811733e-12
+ keta = -0.0962974342888177 lketa = 1.26798662456746e-07 wketa = 5.10577931087838e-08 pketa = -6.90415186675651e-14
+ a1 = 0.0
+ a2 = 2.63306682296493 la2 = -3.65392175475526e-06 wa2 = -8.61068842166555e-07 pa2 = 1.71640124370659e-12
+ ags = 2.81114770247909 lags = -3.00317168385118e-06 wags = -1.27277614170947e-06 pags = 1.65982050580812e-12
+ b0 = -5.25142763609967e-07 lb0 = 1.04042517017215e-12 wb0 = 2.18024251526664e-13 pb0 = -4.54078240025689e-19
+ b1 = 1.09739058232129e-09 lb1 = -4.77784774770859e-14 wb1 = 1.03353572269177e-15 pb1 = 2.57119051808802e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.532927081890699 lvoff = 7.3085599170493e-07 wvoff = 1.08323637791168e-07 pvoff = -3.83020344197045e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -9.72207363067639 lnfactor = 2.32551616713443e-05 wnfactor = 5.62571958286487e-06 pnfactor = -1.08880680984084e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.80670076923077e-05 wcit = -1.08355469408015e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.485738951 leta0 = 9.69238578108438e-07 weta0 = 8.97490964620035e-23 peta0 = 1.73549399148623e-29
+ etab = -0.133215546236516 letab = 2.64546941504003e-07 wetab = 1.77595448696852e-07 petab = -3.54007756514485e-13
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.36833106801906 lpclm = 3.19218178952168e-06 wpclm = 1.37585757763034e-06 ppclm = -1.46627579749537e-12
+ pdiblc1 = 0.375532411367276 lpdiblc1 = 2.8838794189978e-08 wpdiblc1 = 8.37391601679077e-09 ppdiblc1 = -1.66920450050777e-14
+ pdiblc2 = -0.00694737337995754 lpdiblc2 = 7.32822531850026e-09 wpdiblc2 = 4.2558372800508e-09 ppdiblc2 = -4.2274848920911e-15
+ pdiblcb = 1.61421371917477 lpdiblcb = -1.82696087737763e-06 wpdiblcb = -8.63956298715339e-07 ppdiblcb = 8.58200621853297e-13
+ drout = -0.293282617079853 ldrout = 1.70088066536472e-06 wdrout = 3.16124160971165e-07 pdrout = -6.3014230278194e-13
+ pscbe1 = 720796371.089311 lpscbe1 = 157.879603245575 wpscbe1 = 48.2188649321583 ppscbe1 = -9.6116495786139e-5
+ pscbe2 = 1.07385106109966e-08 lpscbe2 = -1.86000686110179e-15 wpscbe2 = -4.15701856385516e-16 ppscbe2 = 4.97246589505542e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.51708125521674e-11 lalpha0 = 1.64070444598945e-16 walpha0 = -1.60477968823172e-17 palpha0 = 1.59408864594873e-23
+ alpha1 = -9.93384736988146e-11 lalpha1 = 1.98010480787033e-16 walpha1 = 2.19543356333498e-21 palpha1 = -2.18080758493604e-27
+ beta0 = -202.001639105538 lbeta0 = 0.000214163831202762 wbeta0 = 0.000120014348768806 pbeta0 = -1.22595061619543e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.93120100905639e-10 lagidl = -2.85212285766503e-15 wagidl = -2.5029874205964e-16 pagidl = 2.04070877929026e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.612971427072123 lkt1 = -8.12183203712924e-09 wkt1 = 8.99248466810301e-08 pkt1 = -2.82589588064781e-14
+ kt2 = -0.0823008217827673 lkt2 = 3.35144258515645e-08 wkt2 = 1.61961184889002e-08 pkt2 = -2.27358070273956e-14
+ at = -285745.954619788 lat = 0.402584132230619 wat = 0.175741811221126 pat = -2.02413490851081e-7
+ ute = -4.80412804441945 lute = 6.56007371686806e-06 wute = 1.8345313272009e-06 pute = -3.00206576383179e-12
+ ua1 = -4.92774614406621e-09 lua1 = 9.94693748164577e-15 wua1 = 2.34711129722896e-15 pua1 = -4.76372523687416e-21
+ ub1 = 4.74651126714728e-18 lub1 = -9.8993281228081e-24 wub1 = -1.93965598315137e-24 pub1 = 4.74618851391443e-30
+ uc1 = 2.19826576922288e-10 luc1 = -3.29578885849329e-16 wuc1 = -7.51402056895185e-17 puc1 = 1.39794341382063e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.104 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.929538946383667 lvth0 = 1.11631718342592e-08 wvth0 = -5.4964212802604e-08 pvth0 = 1.42009964866698e-14
+ k1 = 0.630546320307838 lk1 = -1.89725308634148e-09 wk1 = -1.17911411146093e-07 pk1 = 3.15340709630451e-14
+ k2 = -0.0744147757271736 lk2 = 2.20878737644675e-08 wk2 = 4.78142506842441e-08 pk2 = -1.83184568568631e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1224630.18569422 lvsat = -0.538796170320113 wvsat = -0.565442052593856 pvsat = 2.66244383556583e-7
+ ua = 1.7437277263007e-09 lua = -2.03998849513171e-15 wua = -1.17764438945664e-15 pua = 7.55919510263201e-22
+ ub = -1.31968190557306e-18 lub = 1.62207460798067e-24 wub = 1.17588856953012e-24 pub = -6.10682355138975e-31
+ uc = 7.04290413656642e-11 luc = -2.50022543395987e-17 wuc = -6.43353278308326e-17 puc = 2.20233773020835e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.015596832330387 lu0 = -7.02157589675105e-09 wu0 = -2.18570454592174e-09 pu0 = 2.26672202371729e-15
+ a0 = 3.88213283914244 la0 = -1.58821090686632e-06 wa0 = -1.52640052182606e-06 pa0 = 8.83625889930946e-13
+ keta = -0.0136291570794238 lketa = 4.46811213101213e-08 wketa = 1.43239539183507e-08 pketa = -3.25524003138186e-14
+ a1 = 0.0
+ a2 = -2.86613364592984 la2 = 1.80864304061574e-06 wa2 = 1.72213768433311e-06 pa2 = -8.49595960913526e-13
+ ags = 0.205452758186985 lags = -4.14835879277947e-07 wags = -7.81936461609589e-08 pags = 4.73196318844951e-13
+ b0 = 1.05776915715599e-06 lb0 = -5.31941391377661e-13 wb0 = -5.01565532153337e-13 pb0 = 2.60717636515436e-19
+ b1 = -1.76668707943005e-07 lb1 = 1.28803343299865e-13 wb1 = 9.36586059413534e-14 pb1 = -6.62960968199847e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.543928462211681 lvoff = -3.3882554076264e-07 wvoff = -4.29971325786959e-07 pvoff = 1.51688498333726e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 26.6788220307582 lnfactor = -1.29032312231938e-05 wnfactor = -1.16780628019204e-05 pnfactor = 6.3004364881294e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.58932905741231e-05 lcit = -1.77075241852567e-11 wcit = -2.15267210541638e-11 pcit = 1.06199495114191e-17
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 0.264455062624831 letab = -1.30474385761109e-07 wetab = -3.55197579377524e-07 petab = 1.75235804406859e-13
+ dsub = 0.362722469101819 ldsub = -1.02038132012663e-07 wdsub = -8.38850903282632e-08 pdsub = 8.33262478564963e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.14709555320472 lpclm = -2.9982505955151e-07 wpclm = -2.53232200968339e-07 ppclm = 1.5196098499829e-13
+ pdiblc1 = 1.16248500716365 lpdiblc1 = -7.52871123413203e-07 wpdiblc1 = -3.47988759059294e-07 ppdiblc1 = 3.3729654192965e-13
+ pdiblc2 = 0.00312009841161141 lpdiblc2 = -2.67217697599325e-09 wpdiblc2 = -1.91307069884681e-09 ppdiblc2 = 1.90032582185109e-15
+ pdiblcb = 0.488051315272615 lpdiblcb = -7.08300967410269e-07 wpdiblcb = -4.27646964534492e-07 ppdiblcb = 4.24797980456763e-13
+ drout = 2.07718519040376 ldrout = -6.53795085585443e-07 wdrout = -6.81629508084012e-07 pdrout = 3.60964331329991e-13
+ pscbe1 = 958407257.821378 lpscbe1 = -78.1483197590833 wpscbe1 = -96.4377298643171 ppscbe1 = 4.75763967758022e-5
+ pscbe2 = 4.61851862848446e-08 lpscbe2 = -3.70705367816107e-14 wpscbe2 = -1.75585125069213e-14 ppscbe2 = 1.75258518354874e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 18.9476478061772 lbeta0 = -5.31349155954798e-06 wbeta0 = -7.28230508206667e-06 pbeta0 = 3.85354192337513e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.8544990789564e-09 lagidl = 1.46653248322078e-15 wagidl = 2.86797340045364e-15 pagidl = -1.05678943420959e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.731406532524195 lkt1 = 1.09524258742421e-07 wkt1 = 1.22133617091925e-07 pkt1 = -6.0253154388896e-14
+ kt2 = -0.100048195293156 lkt2 = 5.11435663596272e-08 wkt2 = 3.3583486092534e-08 pkt2 = -4.00073399880541e-14
+ at = 125974.305421817 lat = -0.00639324743858949 wat = -0.0278044992997943 pat = -2.23205850851177e-10
+ ute = 3.48358389471905 lute = -1.6724254853319e-06 wute = -2.24969242817295e-06 pute = 1.05494889288376e-12
+ ua1 = 1.00853785738006e-08 lua1 = -4.96616979935064e-15 wua1 = -5.03818960486036e-15 pua1 = 2.57237479060544e-21
+ ub1 = -1.08912684714139e-17 lub1 = 5.63427272713478e-24 wub1 = 5.66995620747082e-24 pub1 = -2.81272844029384e-30
+ uc1 = -2.46429547484996e-10 luc1 = 1.33571040257153e-16 wuc1 = 1.30309439485697e-16 puc1 = -6.42865982569946e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.105 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.853457644131067 lvth0 = -2.63706256564339e-08 wvth0 = -5.1659753315767e-08 pvth0 = 1.25707810523522e-14
+ k1 = 0.671917546540906 lk1 = -2.23072510937112e-08 wk1 = -1.06544435155784e-07 pk1 = 2.59263097619382e-14
+ k2 = -0.0443411185594837 lk2 = 7.25139588467364e-09 wk2 = 2.10805197888021e-08 pk2 = -5.12969152436754e-15
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 152097.532347528 lvsat = -0.00967505618336287 wvsat = -0.0508386711438604 pvsat = 1.23709805588047e-8
+ ua = -3.21176728642792e-09 lua = 4.04745503457798e-16 wua = 6.9977112982976e-16 pua = -1.70280907190514e-22
+ ub = 2.24513110982347e-18 lub = -1.36583115409023e-25 wub = -1.22287360096497e-25 pub = 2.97571616311615e-32
+ uc = 3.89183171258982e-11 luc = -9.45681666460102e-18 wuc = -3.88627386372953e-17 puc = 9.45678109452218e-24
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00270245356241038 lu0 = 2.00615720702982e-09 wu0 = 4.75372365776541e-09 pu0 = -1.15676160743332e-15
+ a0 = 0.517502082202142 la0 = 7.16893015010951e-08 wa0 = 5.22378037177278e-07 pa0 = -1.27114426810645e-13
+ keta = 0.161533335343541 lketa = -4.17331923768395e-08 wketa = -1.01943398142589e-07 pketa = 2.48067026172214e-14
+ a1 = 0.0
+ a2 = 1.06891451743248 la2 = -1.32665750201105e-7
+ ags = -1.66447624457111 lags = 5.07671155084724e-07 wags = 1.73848168734078e-06 pags = -4.23038656834131e-13
+ b0 = -4.04146836985534e-08 lb0 = 9.83442830183858e-15 wb0 = 5.31052000558932e-14 pb0 = -1.29225131712009e-20
+ b1 = 1.66583825042715e-07 lb1 = -4.05361748182441e-14 wb1 = -8.03629899283572e-14 pb1 = 1.95553692431866e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = 0.128997699621305 lvoff = -1.34124428207829e-07 wvoff = -2.41730782349445e-07 pvoff = 5.88222851153493e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -1.90807716553442 lnfactor = 1.19977245250681e-06 wnfactor = 2.15681736622238e-06 pnfactor = -5.24835624261821e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 2.62181963977308e-05 letab = -2.1588508475031e-11 wetab = 1.33639676417029e-11 petab = -3.2519611579967e-18
+ dsub = -0.30363875647572 ldsub = 2.26703182291309e-07 wdsub = 1.67770180656526e-07 pdsub = -4.08248602205979e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.444148646507052 lpclm = 4.69653615049074e-08 wpclm = 1.08127669747885e-07 ppclm = -2.63115709011107e-14
+ pdiblc1 = -1.16713263793553 lpdiblc1 = 3.96417786384735e-07 wpdiblc1 = 6.62481854051425e-07 ppdiblc1 = -1.61207009401166e-13
+ pdiblc2 = -0.0153041644819908 lpdiblc2 = 6.41721203141068e-09 wpdiblc2 = 3.82614139769362e-09 ppdiblc2 = -9.31045595431972e-16
+ pdiblcb = -1.65110263054523 lpdiblcb = 3.47024961911615e-07 wpdiblcb = 8.55293929068984e-07 ppdiblcb = -2.08125514111788e-13
+ drout = 1.0636610152262 ldrout = -1.53785096051692e-07 wdrout = 9.87623722833648e-08 pdrout = -2.40326381466894e-14
+ pscbe1 = 800069244.26128 lpscbe1 = -0.034160825371373
+ pscbe2 = -6.61067699640808e-08 lpscbe2 = 1.83273523303217e-14 wpscbe2 = 3.54542815693916e-14 ppscbe2 = -8.62737396853262e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.09089376038267 lbeta0 = 5.358957678962e-07 wbeta0 = 1.04361639519408e-06 pbeta0 = -2.53951526373735e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.83748873357367e-09 lagidl = 4.71464633450349e-16 wagidl = 1.43236330889361e-15 pagidl = -3.48548422859554e-22
+ bgidl = 730034204.0064 lbgidl = 133.184385863891
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.506801150159999 lkt1 = -1.28211138236582e-9
+ kt2 = 0.0242671675443682 lkt2 = -1.01859261119115e-08 wkt2 = -9.3757320504542e-08 pkt2 = 2.28147188569342e-14
+ at = 158236.242086396 lat = -0.0223092867488195 wat = -0.0557608877056524 pat = 1.3568742892518e-8
+ ute = 0.364968229524015 lute = -1.33893870295915e-07 wute = -2.19639480984915e-07 pute = 5.34466320239072e-14
+ ua1 = -3.54490332115945e-10 lua1 = 1.8421424695643e-16 wua1 = 3.47377629291368e-16 pua1 = -8.45301775565029e-23
+ ub1 = 6.17482959937584e-19 lub1 = -4.34316865052916e-26 wub1 = -6.20943392504082e-26 pub1 = 1.51099123245158e-32
+ uc1 = 4.743483235632e-11 luc1 = -1.14034251650022e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.106 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.772463663771427 lvth0 = -4.60795388491878e-8
+ k1 = -0.415479539169429 lk1 = 2.4229778094887e-7
+ k2 = 0.438589349394085 lk2 = -1.10263938326212e-07 pk2 = -2.20881053461883e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 92623.7868717143 lvsat = 0.00479716609323078
+ ua = -1.55915274021429e-09 lua = 2.60158501126512e-18
+ ub = 9.27892318000016e-20 lub = 3.87163452505452e-25
+ uc = 6.09622494694279e-15 luc = 1.20053449946548e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0028191509837143 lu0 = 6.62540999984935e-10
+ a0 = -0.39776447742857 la0 = 2.94408435588514e-7
+ keta = -0.184161871607297 lketa = 4.23875878921637e-08 wketa = 1.32348898008484e-23
+ a1 = 0.0
+ a2 = 0.164955374458 la2 = 8.73018597320193e-8
+ ags = -1.62902379023886 lags = 4.99044225752423e-7
+ b0 = 1.23812857142857e-09 lb0 = -3.01283730314285e-16
+ b1 = -1.86798933828571e-10 lb1 = 4.54552789599769e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -0.403685441391143 lvoff = -4.50237804014202e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = -5.59783716277429 lnfactor = 2.09763127071517e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.39713389074943 leta0 = -2.20740146707184e-07 peta0 = 1.0097419586829e-28
+ etab = 0.244655617911143 letab = -5.95492173762617e-08 wetab = 2.98818996284781e-23 petab = 3.10613981430773e-30
+ dsub = 1.53653693089571 ldsub = -2.21081489122281e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.664807054980857 lpclm = -6.72921429629188e-9
+ pdiblc1 = 1.18699067550629 lpdiblc1 = -1.76429872461569e-07 wpdiblc1 = -4.2351647362715e-22
+ pdiblc2 = 0.0300992129326343 lpdiblc2 = -4.63115502190936e-9
+ pdiblcb = -0.782143533009561 lpdiblcb = 1.3557419303548e-7
+ drout = -0.975627884693999 ldrout = 3.42451386277088e-7
+ pscbe1 = 799752699.066858 lpscbe1 = 0.0428666491488912
+ pscbe2 = 2.95389305828885e-08 lpscbe2 = -4.94688114937674e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 11.56376242988 lbeta0 = -5.52523148401942e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.10815918728486e-08 lagidl = 2.72090620315523e-15 wagidl = -2.95822839457879e-31 pagidl = -1.17549435082229e-37
+ bgidl = 1964163557.12 lbgidl = -167.126182664067
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.238369297999999 lkt1 = -6.66017814232761e-8
+ kt2 = 0.235996541485714 lkt2 = -6.17077285080507e-08 wkt2 = -2.64697796016969e-23 pkt2 = 3.15544362088405e-30
+ at = -4339.24200000009 lat = 0.017251506397796
+ ute = -0.316907829714286 lute = 3.20324862070148e-8
+ ua1 = 9.89437705428572e-10 lua1 = -1.42814513843578e-16 wua1 = 3.94430452610506e-31
+ ub1 = 6.03324424e-19 lub1 = -3.99863766873121e-26
+ uc1 = -5.82329727011428e-11 luc1 = 1.43095671820707e-17 wuc1 = -1.23259516440783e-32 puc1 = -2.57139389242375e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.107 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 3.331e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.48711e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__vth0_slope_spectre)
+ vth0 = -0.271654364967343 lvth0 = -1.32888821085291e-07 wvth0 = -3.98278310386429e-07 pvth0 = 6.90367657657628e-14
+ k1 = -3.55748906215231 lk1 = 7.86927427643677e-07 wk1 = 2.03056188465519e-06 pk1 = -3.51973535962361e-13
+ k2 = 0.776126409588245 lk2 = -1.68771937266147e-07 wk2 = -4.41168841059264e-07 pk2 = 7.64713245715306e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 726436.861837209 lvsat = -0.105066724695138 wvsat = -0.291535788567276 pvsat = 5.05342305186745e-8
+ ua = 3.56276519618137e-09 lua = -8.85221426247687e-16 wua = -1.77835174337371e-16 pua = 3.08255934492912e-23
+ ub = 8.79862749666121e-19 lub = 2.50733703065572e-25 wub = -3.2510133643624e-25 pub = 5.63524154551854e-32
+ uc = 8.50235402252939e-13 luc = -1.34316051721212e-19 wuc = -7.01400254704987e-19 puc = 1.21579317350053e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0249695907796761 lu0 = -3.1769719333675e-09 wu0 = -6.3668616419242e-10 pu0 = 1.10361906328787e-16
+ a0 = 8.32068401515669 la0 = -1.21682998921923e-06 wa0 = -2.3328071300386e-06 pa0 = 4.04364122306631e-13
+ keta = 1.11264356092967 lketa = -1.8239807217293e-07 wketa = -3.86463345221317e-07 pketa = 6.69887833339726e-14
+ a1 = 0.0
+ a2 = -4.40683997149522 la2 = 8.7976772140886e-07 wa2 = 2.66744726566008e-06 pa2 = -4.62369974134988e-13
+ ags = -12.5265781191666 lags = 2.3880044980201e-06 wags = 6.47144011416919e-06 pags = -1.12174648650986e-12
+ b0 = -9.43786834473983e-06 lb0 = 1.63585455414051e-12 wb0 = 3.70922238735812e-12 pb0 = -6.42949190179883e-19
+ b1 = -1.58275104845512e-07 lb1 = 2.74481660490793e-14 wb1 = 2.83500848521524e-14 pb1 = -4.9141470081024e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8__voff_slope_spectre)
+ voff = -1.2417827539422 lvoff = 1.40771733922834e-07 wvoff = 5.43094333486554e-07 pvoff = -9.41388855778923e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8__nfactor_slope_spectre)
+ nfactor = 9.86831059126987 lnfactor = -5.83239848675335e-07 wnfactor = -2.25723831182213e-07 pnfactor = 3.91265174494643e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.9160829999519 leta0 = 3.53566242693203e-07 weta0 = 1.06293107742129e-06 peta0 = -1.84246347098052e-13
+ etab = -0.883950891803182 letab = 1.360811778046e-07 wetab = 2.51387450396963e-07 petab = -4.35749978769088e-14
+ dsub = 0.266362313510667 ldsub = -9.11961293991947e-10
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.60108054627701 lpclm = -5.15696988730585e-07 wpclm = -1.76002110450694e-06 ppclm = 3.05078538213025e-13
+ pdiblc1 = 2.54722785653482 lpdiblc1 = -4.12210664946693e-07 wpdiblc1 = -1.45126962854731e-06 ppdiblc1 = 2.51560174873133e-13
+ pdiblc2 = 0.0582974018945875 lpdiblc2 = -9.51897270019641e-09 wpdiblc2 = -3.36595131794213e-08 ppdiblc2 = 5.83447269549454e-15
+ pdiblcb = 1.65062695831742 lpdiblcb = -2.86117378390157e-07 wpdiblcb = -7.75056069871773e-07 ppdiblcb = 1.34346669039433e-13
+ drout = -0.559222936309904 ldrout = 2.70272585334086e-07 wdrout = 9.35131794112962e-07 pdrout = -1.62093874927952e-13
+ pscbe1 = 748810658.381924 lpscbe1 = 8.87305809739428 wpscbe1 = 30.7004083585762 ppscbe1 = -5.32154738405884e-6
+ pscbe2 = -6.16991658561486e-08 lpscbe2 = 1.08681480111731e-14 wpscbe2 = 1.35276716553977e-14 ppscbe2 = -2.34485954940332e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 28.0186167079081 lbeta0 = -3.40477467924677e-06 wbeta0 = -1.00152266064487e-05 pbeta0 = 1.73601934950861e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.56215189917322e-08 lagidl = -3.64113762788948e-15 wagidl = -3.70937252476877e-15 pagidl = 6.4297521469837e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.186819280934522 lkt1 = -7.55373582813718e-08 wkt1 = -2.04704593691399e-07 pkt1 = 3.54830848612796e-14
+ kt2 = -0.12
+ at = 367446.271380506 lat = -0.0471930509205542 wat = -0.0586053616739162 pat = 1.01585361818333e-8
+ ute = -3.56208572623696 lute = 5.94545132434462e-07 wute = 1.67853625105275e-06 pute = -2.90954116684981e-13
+ ua1 = -1.25921172055398e-10 lua1 = 5.05195632617386e-17 wua1 = 2.15887242208684e-16 pua1 = -3.74214627899689e-23
+ ub1 = 3.7264e-19
+ uc1 = 2.53798686275156e-10 luc1 = -3.97773765215631e-17 wuc1 = -1.38499172747403e-16 puc1 = 2.40071696056894e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 5.24898e-11
+ cgso = 5.24898e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 9.5483718e-12
+ cgdl = 9.5483718e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.4325e-8
+ dwc = -3.2175e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006679036719
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 8.9499956e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.0 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4181113
+ k1 = 0.47213
+ k2 = -0.0321739
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161140.0
+ ua = -1.3019497e-9
+ ub = 2.64393e-18
+ uc = 7.0152e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03208538
+ a0 = 1.9632567
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5148757
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11559919
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.1534679
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0047977
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.4345657e-5
+ alpha1 = 0.0
+ beta0 = 17.822982
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25364
+ kt2 = -0.034423
+ at = 333080.0
+ ute = -1.0777
+ ua1 = 2.6823e-9
+ ub1 = -2.4433e-18
+ uc1 = -1.9223e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.1 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.039508629e-01 lvth0 = 1.134335973e-07 wvth0 = 9.747549271e-08 pvth0 = -7.808371819e-13
+ k1 = 5.494703645e-01 lk1 = -6.195427239e-07 wk1 = -5.323840001e-07 pk1 = 4.264715271e-12
+ k2 = -5.912813589e-02 lk2 = 2.159196020e-07 wk2 = 1.855435259e-07 pk2 = -1.486314969e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.304176524e+04 lvsat = 7.057197193e-01 wvsat = 6.064374137e-01 pvsat = -4.857927546e-6
+ ua = -1.340324789e-09 lua = 3.074074899e-16 wua = 2.641606831e-16 pua = -2.116085568e-21
+ ub = 2.675649026e-18 lub = -2.540884285e-25 wub = -2.183426723e-25 pub = 1.749055811e-30
+ uc = 6.984078634e-11 luc = 2.493008176e-18 wuc = 2.142285938e-18 puc = -1.716099573e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.162412689e-02 lu0 = 3.694914159e-09 wu0 = 3.175104968e-09 pu0 = -2.543449585e-14
+ a0 = 2.000299418e+00 la0 = -2.967343957e-07 wa0 = -2.549891048e-07 pa0 = 2.042615723e-12
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.008643009e-01 lags = 1.122397138e-07 wags = 9.644956754e-08 pags = -7.726189057e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.120409948e-01 lvoff = -2.850327846e-08 wvoff = -2.449337038e-08 pvoff = 1.962065928e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.261889959e+00 lnfactor = -8.685257477e-07 wnfactor = -7.463395080e-07 pnfactor = 5.978627263e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.416657520e-01 lpclm = -1.134827673e-06 wpclm = -9.751774541e-07 ppclm = 7.811756514e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.870867443e-03 lpdiblc2 = 1.543508488e-08 wpdiblc2 = 1.326364093e-08 ppdiblc2 = -1.062497220e-13
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.387872744e-04 lalpha0 = -4.361100204e-10 walpha0 = -3.747570396e-10 palpha0 = 3.002028742e-15
+ alpha1 = 0.0
+ beta0 = 1.812625487e+01 lbeta0 = -2.429397649e-06 wbeta0 = -2.087624289e-06 pbeta0 = 1.672312313e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.532200231e-01 lkt1 = -3.364267089e-09 wkt1 = -2.890974103e-09 pkt1 = 2.315843715e-14
+ kt2 = -3.413547734e-02 lkt2 = -2.303229007e-09 wkt2 = -1.979205347e-09 pkt2 = 1.585462235e-14
+ at = 6.184327776e+05 lat = -2.285846960e+00 wat = -1.964268648e+00 pat = 1.573497043e-5
+ ute = -9.493378244e-01 lute = -1.028258044e-06 wute = -8.836002898e-07 pute = 7.078168482e-12
+ ua1 = 2.420622075e-09 lua1 = 2.096197186e-15 wua1 = 1.801299249e-15 pua1 = -1.442948776e-20
+ ub1 = -1.549718345e-18 lub1 = -7.158125206e-24 wub1 = -6.151103360e-24 pub1 = 4.927402857e-29
+ uc1 = -1.087192054e-11 luc1 = -6.689715711e-17 wuc1 = -5.748590812e-17 puc1 = 4.604966156e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.2 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.321459564e-01 lvth0 = 3.543554001e-10 wvth0 = -1.949509854e-07 pvth0 = 3.919684513e-13
+ k1 = 3.594104930e-01 lk1 = 1.427113968e-07 wk1 = 1.064768000e-06 pk1 = -2.140822541e-12
+ k2 = 6.612547593e-03 lk2 = -4.773998315e-08 wk2 = -3.710870518e-07 pk2 = 7.461076263e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.535984092e+05 lvsat = -8.205407570e-01 wvsat = -1.212874827e+00 pvsat = 2.438606128e-6
+ ua = -1.302525680e-09 lua = 1.558103804e-16 wua = -5.283213661e-16 pua = 1.062242939e-21
+ ub = 2.594422390e-18 lub = 7.167911566e-26 wub = 4.366853446e-25 pub = -8.779995538e-31
+ uc = 6.796662443e-11 luc = 1.000952193e-17 wuc = -4.284571875e-18 puc = 8.614560212e-24
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.076770586e-02 lu0 = 7.129676352e-09 wu0 = -6.350209935e-09 pu0 = 1.276773210e-14
+ a0 = 1.900878686e+00 la0 = 1.020023895e-07 wa0 = 5.099782096e-07 pa0 = -1.025362188e-12
+ keta = 1.855080090e-01 lketa = -7.439984209e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.747436646e-01 lags = 3.623953020e-06 wags = -1.928991351e-07 pags = 3.878430010e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.224166343e-01 lvoff = 1.310926146e-08 wvoff = 4.898674077e-08 pvoff = -9.849274098e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 7.073644128e-01 lnfactor = 1.355454409e-06 wnfactor = 1.492679016e-06 pnfactor = -3.001180430e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 8.384947203e-01 ldsub = -1.116930925e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.135910341e-01 lpclm = 6.910251931e-07 wpclm = 1.950354908e-06 ppclm = -3.921383578e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 4.736927973e-03 lpdiblc2 = 7.951062517e-09 wpdiblc2 = -2.652728186e-08 ppdiblc2 = 5.333575290e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.619115086e-05 lalpha0 = 3.859764520e-10 walpha0 = 7.495140793e-10 palpha0 = -1.506973008e-15
+ alpha1 = 0.0
+ beta0 = 1.372440306e+01 lbeta0 = 1.522466922e-05 wbeta0 = 4.175248578e-06 pbeta0 = -8.394754790e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.544900068e-01 lkt1 = 1.729129739e-09 wkt1 = 5.781948205e-09 pkt1 = -1.162518506e-14
+ kt2 = -3.979131572e-02 lkt2 = 2.038007638e-08 wkt2 = 3.958410694e-09 pkt2 = -7.958780542e-15
+ at = 4.556946537e+04 lat = 1.167863972e-02 wat = 3.928537295e+00 pat = -7.898717086e-6
+ ute = -1.242439401e+00 lute = 1.472551399e-07 wute = 1.767200580e-06 pute = -3.553133485e-12
+ ua1 = 2.632835910e-09 lua1 = 1.245092379e-15 wua1 = -3.602598497e-15 pua1 = 7.243384538e-21
+ ub1 = -2.899948760e-18 lub1 = -1.742891103e-24 wub1 = 1.230220672e-23 pub1 = -2.473481683e-29
+ uc1 = -2.031787642e-11 luc1 = -2.901320647e-17 wuc1 = 1.149718162e-16 puc1 = -2.311623337e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.3 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.296412904e-01 lvth0 = 5.390236789e-9
+ k1 = 4.289650540e-01 lk1 = 2.864996428e-9
+ k2 = -1.322128542e-02 lk2 = -7.862078495e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.825027700e+04 lvsat = 5.477019766e-2
+ ua = -9.408298839e-10 lua = -5.714151863e-16
+ ub = 2.567681588e-18 lub = 1.254441734e-25
+ uc = 5.919376580e-11 luc = 2.764823148e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.856590003e-02 lu0 = -8.549372850e-9
+ a0 = 2.194610781e+00 la0 = -4.885753589e-7
+ keta = -1.435097460e-01 lketa = -8.247532269e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.402628058e-01 lags = 1.382121011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.171097954e-01 lvoff = 2.439331107e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 9.970702915e-01 lnfactor = 7.729717692e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.944506760e-04 leta0 = -1.899025292e-10
+ etab = -5.430717720e-04 letab = 8.660010478e-11
+ dsub = -6.340633544e-02 ldsub = 6.964313374e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.292005660e-01 lpclm = 1.808402000e-9
+ pdiblc1 = 0.39
+ pdiblc2 = 6.955794500e-03 lpdiblc2 = 3.489809478e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.887537269e-04 lalpha0 = -1.266157192e-10
+ alpha1 = 0.0
+ beta0 = 2.119341263e+01 lbeta0 = 2.074785711e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.505779880e-01 lkt1 = -6.136375327e-9
+ kt2 = -4.652898820e-02 lkt2 = 3.392684067e-8
+ at = 3.027262960e+04 lat = 4.243445773e-2
+ ute = -1.329885400e+00 lute = 3.230740652e-7
+ ua1 = 3.274737440e-09 lua1 = -4.551483686e-17
+ ub1 = -3.913337000e-18 lub1 = 2.946272922e-25
+ uc1 = 1.290785360e-11 luc1 = -9.581685925e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.4 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.400250589e-01 lvth0 = -5.103599606e-9
+ k1 = 4.339445200e-01 lk1 = -2.167251912e-9
+ k2 = -1.418804385e-02 lk2 = -6.885072422e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.026880832e+04 lvsat = 6.283626991e-2
+ ua = -1.198824854e-09 lua = -3.106854690e-16
+ ub = 2.616425016e-18 lub = 7.618406483e-26
+ uc = 1.089428312e-10 luc = -2.262817401e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.375954300e-02 lu0 = -3.692068436e-9
+ a0 = 1.969380632e+00 la0 = -2.609577707e-7
+ keta = -4.454529355e-01 lketa = 2.226684646e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.902775804e+00 lags = -8.033146257e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.149895327e-01 lvoff = 2.965935843e-10
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.194371862e+00 lnfactor = 5.735788021e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 8.114866480e-04 leta0 = -4.092390825e-10
+ etab = -8.606660737e-04 letab = 4.075609060e-10
+ dsub = 2.435057895e-01 ldsub = 3.862659439e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.109362400e-02 lpclm = 2.951797104e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.029564680e-02 lpdiblc2 = 1.145547439e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.483090005e-05 lalpha0 = 9.933890479e-11
+ alpha1 = 0.0
+ beta0 = 1.835426046e+01 lbeta0 = 3.076725761e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.502470760e-01 lkt1 = -6.470794994e-9
+ kt2 = -4.901692000e-04 lkt2 = -1.259998981e-8
+ at = 7.237126840e+04 lat = -1.104266450e-4
+ ute = -1.004685520e+00 lute = -5.572933488e-9
+ ua1 = 4.088120720e-09 lua1 = -8.675199796e-16
+ ub1 = -4.763807960e-18 lub1 = 1.154113244e-24
+ uc1 = -1.743066693e-10 luc1 = 9.338213757e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.5 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.053773090e-01 lvth0 = -3.847245853e-8
+ k1 = 2.731315200e-01 lk1 = 7.994386589e-8
+ k2 = 2.685855531e-02 lk2 = -2.784346596e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.935343216e+04 lvsat = 3.266766098e-2
+ ua = -1.672033646e-09 lua = -6.906505991e-17
+ ub = 2.983232042e-18 lub = -1.111076028e-25
+ uc = 7.538546830e-11 luc = -5.493784512e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.311010088e-02 lu0 = -3.360463289e-9
+ a0 = 1.296832240e+00 la0 = 8.244543826e-8
+ keta = -1.428146283e-02 lketa = 2.512310660e-9
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.715370800e+00 lags = -7.076256305e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.192914701e-01 lvoff = 2.493162827e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.795148014e+00 lnfactor = 2.668224990e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -5.996306819e-03 leta0 = 3.066820262e-09 weta0 = -1.525114254e-24 peta0 = -4.252453317e-31
+ etab = 2.833070331e-02 letab = -1.449755230e-08 wetab = 5.169878828e-24 petab = 5.472722530e-30
+ dsub = 1.760787113e+00 ldsub = -3.884579000e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.596832880e-01 lpclm = -7.284898085e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 6.953949600e-03 lpdiblc2 = 1.820825334e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.658135538e-03 lalpha0 = 1.438798253e-09 walpha0 = -4.135903063e-25 palpha0 = 3.944304526e-31
+ alpha1 = 0.0
+ beta0 = 1.719950301e+01 lbeta0 = 3.666344913e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.525689680e-01 lkt1 = -5.285236939e-9
+ kt2 = -2.883937520e-02 lkt2 = 1.875114777e-9
+ at = 8.981221360e+04 lat = -9.015773264e-3
+ ute = -3.364764000e-01 lute = -3.467605102e-7
+ ua1 = 4.368482088e-09 lua1 = -1.010672494e-15
+ ub1 = -4.381560808e-18 lub1 = 9.589378486e-25
+ uc1 = 5.561182016e-11 luc1 = -2.401424313e-17 wuc1 = -2.465190329e-32 puc1 = 5.877471754e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.6 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 6.162803797e-01 lvth0 = -6.737379875e-8
+ k1 = 2.569146857e-01 lk1 = 8.416997290e-8
+ k2 = 3.072747161e-02 lk2 = -2.885170554e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.954686771e+05 lvsat = -1.979718634e-4
+ ua = -6.981024429e-10 lua = -3.228715315e-16
+ ub = 1.429150534e-18 lub = 2.938860382e-25
+ uc = 8.960922466e-11 luc = -9.200495420e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.561932686e-02 lu0 = -1.408367579e-9
+ a0 = 6.005713143e+00 la0 = -1.144688925e-6
+ keta = 3.021383089e-01 lketa = -7.994668186e-08 wketa = 1.588186776e-22 pketa = -3.155443621e-29
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.277775429e+00 lags = 8.541882767e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.759880884e-01 lvoff = 1.726830156e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.114708772e+00 lnfactor = 1.835449655e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.893770899e-01 leta0 = 5.085585235e-08 peta0 = 6.310887242e-30
+ etab = -6.126409553e-02 letab = 8.850852274e-9
+ dsub = 1.292577563e-01 ldsub = 3.671865043e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.011325514e+00 lpclm = -1.644869450e-7
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 1.457542571e-02 lpdiblc2 = -1.653313411e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.906043181e-03 lalpha0 = -1.574826721e-9
+ alpha1 = 0.0
+ beta0 = 3.744754421e+01 lbeta0 = -1.610294622e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.620297143e-01 lkt1 = -2.887976646e-8
+ kt2 = -3.810094857e-02 lkt2 = 4.288680798e-9
+ at = -1.210119714e+04 lat = 1.754286158e-2
+ ute = -1.022327429e+00 lute = -1.680277321e-7
+ ua1 = 1.775331440e-09 lua1 = -3.348974353e-16
+ ub1 = -2.283428800e-18 lub1 = 4.121646473e-25
+ uc1 = -1.411542557e-10 luc1 = 2.726299624e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.7 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 1.128974073e-01 lvth0 = 2.857099578e-8
+ k1 = 1.097236267e+00 lk1 = -7.599532043e-8
+ k2 = -2.061792656e-01 lk2 = 1.630271857e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.276902600e+05 lvsat = -6.339405556e-3
+ ua = -3.793134041e-09 lua = 2.670414910e-16
+ ub = 5.948734600e-18 lub = -5.675466848e-25
+ uc = 2.262694353e-10 luc = -3.524793157e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.199305800e-02 lu0 = -7.172007348e-10
+ a0 = 0.0
+ keta = 2.323739224e-01 lketa = -6.664958979e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.505873333e-01 lags = 4.826233427e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.286910051e-01 lvoff = 8.253477489e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -2.225938087e-01 lnfactor = 6.290348373e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 6.493980999e-02 leta0 = 2.383051218e-9
+ etab = -9.420281110e-02 letab = 1.512897146e-8
+ dsub = 6.533059590e-01 ldsub = -6.316493702e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.990366667e-02 lpclm = 1.494805913e-8
+ pdiblc1 = 4.294484535e+00 lpdiblc1 = -6.279287523e-7
+ pdiblc2 = 7.877401933e-02 lpdiblc2 = -1.240158328e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.974575979e-03 lalpha0 = -2.536890724e-10
+ alpha1 = 0.0
+ beta0 = 3.185758335e+01 lbeta0 = -5.448480825e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.900488667e-01 lkt1 = -4.479316013e-9
+ kt2 = 3.135944000e-02 lkt2 = -8.950469264e-9
+ at = 5.954280000e+04 lat = 3.887515720e-3
+ ute = -3.099299333e+00 lute = 2.278431129e-7
+ ua1 = -3.102292360e-09 lua1 = 5.947776610e-16 wua1 = -6.902532921e-31 pua1 = 1.410593221e-37
+ ub1 = 3.150130800e-18 lub1 = -6.234718125e-25 wub1 = -1.469367939e-39 pub1 = -1.751623080e-46
+ uc1 = 6.131370000e-12 luc1 = -8.096440220e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.8 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.848415475e-01 wvth0 = 2.290173319e-7
+ k1 = 6.538401246e-01 wk1 = -1.250828899e-6
+ k2 = -9.550250718e-02 wk2 = 4.359319668e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.584559308e+04 wvsat = 1.424816378e+0
+ ua = -1.392111445e-09 wua = 6.206418982e-16
+ ub = 2.718453416e-18 wub = -5.129931110e-25
+ uc = 6.942080777e-11 wuc = 5.033271399e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.100167215e-02 wu0 = 7.459865531e-9
+ a0 = 2.050288057e+00 wa0 = -5.990934010e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.819561101e-01 wags = 2.266069348e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.072392592e-01 wvoff = -5.754683745e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.408204040e+00 wnfactor = -1.753514428e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.328417395e-01 wpclm = -2.291166040e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.706333615e-04 wpdiblc2 = 3.116274227e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.122554897e-04 walpha0 = -8.804865197e-10
+ alpha1 = 0.0
+ beta0 = 1.853551744e+01 wbeta0 = -4.904844606e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.526532700e-01 wkt1 = -6.792303964e-9
+ kt2 = -3.374746946e-02 wkt2 = -4.650115791e-9
+ at = 1.003512433e+06 wat = -4.615022221e+0
+ ute = -7.761148308e-01 wute = -2.076006750e-6
+ ua1 = 2.067491308e-09 wua1 = 4.232127855e-15
+ ub1 = -3.438421692e-19 wub1 = -1.445193290e-23
+ uc1 = 3.977465385e-13 wuc1 = -1.350623519e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.9 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.848415475e-01 wvth0 = 2.290173319e-7
+ k1 = 6.538401246e-01 wk1 = -1.250828899e-6
+ k2 = -9.550250718e-02 wk2 = 4.359319668e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.584559308e+04 wvsat = 1.424816378e+0
+ ua = -1.392111445e-09 wua = 6.206418982e-16
+ ub = 2.718453416e-18 wub = -5.129931110e-25
+ uc = 6.942080777e-11 wuc = 5.033271399e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.100167215e-02 wu0 = 7.459865531e-9
+ a0 = 2.050288057e+00 wa0 = -5.990934010e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.819561101e-01 wags = 2.266069348e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.072392592e-01 wvoff = -5.754683745e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.408204040e+00 wnfactor = -1.753514428e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.328417395e-01 wpclm = -2.291166040e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.706333615e-04 wpdiblc2 = 3.116274227e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.122554897e-04 walpha0 = -8.804865197e-10
+ alpha1 = 0.0
+ beta0 = 1.853551744e+01 wbeta0 = -4.904844606e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.526532700e-01 wkt1 = -6.792303964e-9
+ kt2 = -3.374746946e-02 wkt2 = -4.650115791e-9
+ at = 1.003512433e+06 wat = -4.615022221e+0
+ ute = -7.761148308e-01 wute = -2.076006750e-6
+ ua1 = 2.067491308e-09 wua1 = 4.232127855e-15
+ ub1 = -3.438421692e-19 wub1 = -1.445193290e-23
+ uc1 = 3.977465385e-13 wuc1 = -1.350623519e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.10 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.186186106e-01 lvth0 = 2.655937107e-07 wvth0 = 5.865315285e-07 pvth0 = -1.433846437e-12
+ k1 = 1.043546798e+00 lk1 = -1.562957583e-06 wk1 = -3.644586874e-06 pk1 = 9.600405734e-12
+ k2 = -2.374048848e-01 lk2 = 5.691136756e-07 wk2 = 1.308643546e-06 pk2 = -3.500097061e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.297178753e+05 lvsat = 3.363781751e-01 wvsat = 2.802470315e+00 pvsat = -5.525218879e-6
+ ua = -1.629846028e-09 lua = 9.534583169e-16 wua = 1.724837350e-15 pua = -4.428486280e-21
+ ub = 2.613463154e-18 lub = 4.210739420e-25 wub = 3.056153890e-25 pub = -3.283111250e-30
+ uc = 1.253293868e-10 luc = -2.242269471e-16 wuc = -3.991497512e-16 puc = 1.621016430e-21
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.396846984e-02 lu0 = 2.820736117e-08 wu0 = 4.045335105e-08 pu0 = -1.323236730e-13
+ a0 = 2.043295005e+00 la0 = 2.804633571e-08 wa0 = -4.703658793e-07 pa0 = -5.162745983e-13
+ keta = 1.054644942e-01 lketa = -4.229759003e-07 wketa = 5.509915409e-07 pketa = -2.209806674e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.179047199e-01 lags = 4.411101845e-06 wags = 1.480936464e-06 pags = -5.030614009e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -8.697351308e-02 lvoff = -8.127780151e-08 wvoff = -1.949913009e-07 pvoff = 5.512347650e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.163203045e+00 lnfactor = -3.027999010e-06 wnfactor = -8.528804583e-06 pnfactor = 2.717297870e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.717431654e-06 lcit = 5.100453139e-11 wcit = 8.754234840e-11 pcit = -3.510973425e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 1.190469989e+00 ldsub = -2.528562939e-06 wdsub = -2.422874560e-06 pdsub = 9.717180710e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.773409426e-01 lpclm = 6.236514962e-07 wpclm = -1.429048993e-06 ppclm = -3.457606629e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -7.961117476e-03 lpdiblc2 = 3.301425991e-08 wpdiblc2 = 6.088161870e-08 ppdiblc2 = -1.191905258e-13
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.076305106e-04 lalpha0 = -3.825110588e-10 walpha0 = -1.823743400e-09 palpha0 = 3.783026046e-15
+ alpha1 = 0.0
+ beta0 = 1.581270064e+01 lbeta0 = 1.092012908e-05 wbeta0 = -1.019986106e-05 pbeta0 = 2.123619298e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.795734084e-01 lkt1 = 1.079659070e-07 wkt1 = 1.784473053e-07 pkt1 = -7.429219767e-13
+ kt2 = -1.800463123e-02 lkt2 = -6.313822702e-08 wkt2 = -1.460135000e-07 pkt2 = 5.669519887e-13
+ at = 1.978121148e+06 lat = -3.908765710e+00 wat = -9.374472093e+00 pat = 1.908824966e-5
+ ute = -5.442381326e-01 lute = -9.299646858e-07 wute = -3.038972583e-06 pute = 3.862070768e-12
+ ua1 = -7.067160516e-10 lua1 = 1.112623604e-14 wua1 = 1.938570836e-14 pua1 = -6.077494999e-20
+ ub1 = 5.364266705e-18 lub1 = -2.289294145e-23 wub1 = -4.458576006e-23 pub1 = 1.208547272e-28
+ uc1 = 2.364566198e-11 luc1 = -9.323808965e-17 wuc1 = -1.876577948e-16 puc1 = 2.109392834e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.11 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.697118313e-01 lvth0 = -3.819431880e-08 wvth0 = -2.758315786e-07 pvth0 = 3.000208261e-13
+ k1 = 1.085111631e-01 lk1 = 3.170250637e-07 wk1 = 2.205892426e-06 pk1 = -2.162567947e-12
+ k2 = 1.046061518e-01 lk2 = -1.185337146e-07 wk2 = -8.110828382e-07 pk2 = 7.618248076e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.306448244e+03 lvsat = 6.288767019e-02 wvsat = 8.221713681e-02 pvsat = -5.587783977e-8
+ ua = -8.695680040e-10 lua = -5.751566780e-16 wua = -4.905418394e-16 pua = 2.575511907e-23
+ ub = 2.878397213e-18 lub = -1.116024753e-25 wub = -2.138857611e-24 pub = 1.631746163e-30
+ uc = -8.624971096e-11 luc = 2.011739869e-16 wuc = 1.001181989e-15 puc = -1.194490566e-21
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.466544444e-02 lu0 = -1.340597595e-08 wu0 = -4.198712889e-08 pu0 = 3.343115594e-14
+ a0 = 2.528528788e+00 la0 = -9.475647080e-07 wa0 = -2.298574688e-06 pa0 = 3.159522033e-12
+ keta = 1.597890140e-01 lketa = -5.322007798e-07 wketa = -2.087802509e-06 pketa = 3.095752643e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.776907494e-01 lags = 1.605117594e-06 wags = -2.576408636e-07 pags = -1.535030434e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.424255136e-01 lvoff = 3.021399080e-08 wvoff = 1.742645438e-07 pvoff = -1.911910362e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -4.667114723e-01 lnfactor = 2.259707118e-06 wnfactor = 1.007616134e-05 pnfactor = -1.023416578e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.048786331e-05 lcit = -3.586403466e-11 wcit = -1.750846968e-10 pcit = 1.769405946e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 7.633336395e-04 leta0 = -5.294586156e-10 weta0 = -1.162531212e-09 peta0 = 2.337385255e-15
+ etab = -5.914993773e-04 letab = 1.839686480e-10 wetab = 3.333586851e-10 petab = -6.702509723e-16
+ dsub = 1.896373989e-01 ldsub = -5.162889328e-07 wdsub = -1.741864502e-06 pdsub = 8.347941888e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.257307081e+00 lpclm = -1.145608421e-06 wpclm = -7.077125410e-06 ppclm = 7.898415814e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.062535902e-02 lpdiblc2 = -4.355709728e-09 wpdiblc2 = -2.525999779e-08 ppdiblc2 = 5.400580828e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.625105526e-04 lalpha0 = -9.073287141e-11 walpha0 = 1.806488263e-10 palpha0 = -2.470049650e-16
+ alpha1 = 0.0
+ beta0 = 2.066982985e+01 lbeta0 = 1.154385083e-06 wbeta0 = 3.604160624e-06 pbeta0 = -6.518173012e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.146409778e-01 lkt1 = -2.258723796e-08 wkt1 = -2.473778003e-07 pkt1 = 1.132419805e-13
+ kt2 = -1.442129240e-01 lkt2 = 1.906161663e-07 wkt2 = 6.724220243e-07 pkt2 = -1.078594477e-12
+ at = -7.658617393e+02 lat = 6.998451174e-02 wat = 2.136581109e-01 pat = -1.896449293e-7
+ ute = -1.419053002e+00 lute = 8.289380911e-07 wute = 6.137985649e-07 pute = -3.482190902e-12
+ ua1 = 3.748199640e-09 lua1 = 2.169182545e-15 wua1 = -3.259148076e-15 pua1 = -1.524520163e-20
+ ub1 = -4.708151405e-18 lub1 = -2.641337598e-24 wub1 = 5.471224181e-24 pub1 = 2.021015471e-29
+ uc1 = 1.746472790e-10 luc1 = -3.968419409e-16 wuc1 = -1.113357596e-15 puc1 = 2.072151303e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.12 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.333120577e-01 lvth0 = -1.408707601e-09 wvth0 = 4.620995066e-08 pvth0 = -2.543434335e-14
+ k1 = 4.514845313e-01 lk1 = -2.958382216e-08 wk1 = -1.207392986e-07 pk1 = 1.887260738e-13
+ k2 = -8.231423878e-03 lk2 = -4.500060587e-09 wk2 = -4.100328710e-08 pk2 = -1.641758671e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.816690595e+05 lvsat = -1.143337848e-01 wvsat = -1.179859339e+00 pvsat = 1.219576647e-6
+ ua = -5.836471811e-10 lua = -8.641082616e-16 wua = -4.234667791e-15 pua = 3.809568806e-21
+ ub = 2.215394090e-18 lub = 5.584284799e-25 wub = 2.760556531e-24 pub = -3.319601768e-30
+ uc = 1.393033384e-10 luc = -2.676992478e-17 wuc = -2.089911051e-16 puc = 2.851036267e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.021542765e-02 lu0 = -8.908788978e-09 wu0 = -4.444005034e-08 pu0 = 3.591007836e-14
+ a0 = 2.002257724e+00 la0 = -4.157151709e-07 wa0 = -2.263143920e-07 pa0 = 1.065295778e-12
+ keta = -7.076898512e-01 lketa = 3.444733613e-07 wketa = 1.805147145e-06 pketa = -8.384622771e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.237255728e-01 lags = 2.266014802e-06 wags = 1.913000913e-05 pags = -2.112818951e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.108157119e-01 lvoff = -1.730874841e-09 wvoff = -2.873112141e-08 pvoff = 1.395638302e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 6.156082103e-01 lnfactor = 1.165914847e-06 wnfactor = 3.984006410e-06 pnfactor = -4.077434013e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.478836202e-04 leta0 = -2.106647808e-10 weta0 = 2.502916291e-09 peta0 = -1.366915991e-15
+ etab = -7.654270721e-04 letab = 3.597399764e-10 wetab = -6.555919528e-10 petab = 3.291825424e-16
+ dsub = -1.670482755e+00 ldsub = 1.363548495e-06 wdsub = 1.317522724e-05 pdsub = -6.727271031e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.198471667e-01 lpclm = 7.514436613e-07 wpclm = 3.846263824e-06 ppclm = -3.140761346e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.901748210e-04 lpdiblc2 = 5.987967421e-09 wpdiblc2 = 6.818580219e-08 ppdiblc2 = -4.043051717e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.196680708e-04 lalpha0 = 1.944368455e-10 walpha0 = 5.839893905e-10 palpha0 = -6.546209392e-16
+ alpha1 = 0.0
+ beta0 = 1.805258342e+01 lbeta0 = 3.799374330e-06 wbeta0 = 2.076639166e-06 pbeta0 = -4.974459826e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.173339226e-01 lkt1 = -1.986574789e-08 wkt1 = -2.265626281e-07 pkt1 = 9.220616747e-14
+ kt2 = 9.152968183e-02 lkt2 = -4.762531107e-08 wkt2 = -6.334324475e-07 pkt2 = 2.411020527e-13
+ at = 8.178866141e+03 lat = 6.094496974e-02 wat = 4.418780298e-01 pat = -4.202839793e-7
+ ute = -2.481107479e-01 lute = -3.544161511e-07 wute = -5.207995930e-06 pute = 2.401314615e-12
+ ua1 = 9.514008115e-09 lua1 = -3.657743500e-15 wua1 = -3.734990977e-14 pua1 = 1.920692214e-20
+ ub1 = -1.237295257e-17 lub1 = 5.104710462e-24 wub1 = 5.237868831e-23 pub1 = -2.719452853e-29
+ uc1 = -5.389396767e-10 luc1 = 3.243090365e-16 wuc1 = 2.510006001e-15 puc1 = -1.589619948e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.13 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.331111927e-01 lvth0 = -5.236614593e-08 wvth0 = -1.909103482e-07 pvth0 = 9.563928123e-14
+ k1 = 2.555436801e-01 lk1 = 7.046357643e-08 wk1 = 1.210685338e-07 pk1 = 6.525899454e-14
+ k2 = 3.010826017e-02 lk2 = -2.407630326e-08 wk2 = -2.236983086e-08 pk2 = -2.593182947e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.297686431e+05 lvsat = 1.468063062e-01 wvsat = 2.747416673e+00 pvsat = -7.856904850e-7
+ ua = -1.912290361e-09 lua = -1.857030541e-16 wua = 1.653843131e-15 pua = 8.028951290e-22
+ ub = 2.990337962e-18 lub = 1.627421392e-25 wub = -4.891466205e-26 pub = -1.885085777e-30
+ uc = 1.412058887e-10 luc = -2.774136697e-17 wuc = -4.530847367e-16 puc = 1.531445710e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.893639592e-02 lu0 = -3.149715377e-09 wu0 = 2.873032417e-08 pu0 = -1.450714864e-15
+ a0 = 3.047767317e-01 la0 = 4.510186236e-07 wa0 = 6.828962900e-06 pa0 = -2.537128807e-12
+ keta = -1.437341228e-01 lketa = 5.651756640e-08 wketa = 8.911068031e-07 pketa = -3.717532787e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.316756318e+00 lags = -2.427946696e-06 wags = -4.544162742e-05 pags = 1.184208811e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.244823715e-01 lvoff = 5.247321578e-09 wvoff = 3.573234884e-08 pvoff = -1.895866489e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 3.239326621e+00 lnfactor = -1.737557741e-07 wnfactor = -9.941220074e-06 pnfactor = 3.032786630e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.171196991e-02 leta0 = 5.998157005e-09 weta0 = 3.934463227e-08 peta0 = -2.017829617e-14
+ etab = -4.800475600e-02 letab = 2.448014133e-08 wetab = 5.254665845e-07 petab = -2.683088007e-13
+ dsub = 1.943666626e+00 ldsub = -4.818361791e-07 wdsub = -1.258878557e-06 pdsub = 6.427833910e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.376085782e+00 lpclm = -2.676797023e-07 wpclm = -4.931464028e-06 ppclm = 1.341146496e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.278808272e-02 lpdiblc2 = -3.424043515e-10 wpdiblc2 = -4.016013044e-08 ppdiblc2 = 1.489091603e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.138920428e-03 lalpha0 = 2.757267099e-09 walpha0 = 1.707685491e-08 palpha0 = -9.075878072e-15
+ alpha1 = 0.0
+ beta0 = 1.743969906e+01 lbeta0 = 4.112313081e-06 wbeta0 = -1.653425558e-06 pbeta0 = -3.069888778e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.672173493e-01 lkt1 = -4.545527026e-08 wkt1 = -5.875306704e-07 pkt1 = 2.765164499e-13
+ kt2 = 7.667981142e-03 lkt2 = -4.805526701e-09 wkt2 = -2.513038635e-07 pkt2 = 4.598719771e-14
+ at = 1.856314811e+05 lat = -2.966233548e-02 wat = -6.595863010e-01 pat = 1.421237080e-7
+ ute = 1.996209953e+00 lute = -1.500366301e-06 wute = -1.605739642e-05 pute = 7.941018503e-12
+ ua1 = 9.687473754e-09 lua1 = -3.746315055e-15 wua1 = -3.661407698e-14 pua1 = 1.883120591e-20
+ ub1 = -8.512256103e-18 lub1 = 3.133438844e-24 wub1 = 2.843426067e-23 pub1 = -1.496850378e-29
+ uc1 = 3.309565358e-10 luc1 = -1.198599696e-16 wuc1 = -1.895376652e-15 puc1 = 6.597684348e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.14 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 6.621173163e-01 lvth0 = -8.598514176e-08 wvth0 = -3.155254289e-07 pvth0 = 1.281139713e-13
+ k1 = 9.113905785e-02 lk1 = 1.133074210e-07 wk1 = 1.141141401e-06 pk1 = -2.005719946e-13
+ k2 = 4.644887520e-02 lk2 = -2.833466754e-08 wk2 = -1.082206399e-07 pk2 = -3.559108644e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.024081324e+05 lvsat = -1.793896152e-02 wvsat = -7.361337813e-01 pvsat = 1.221227634e-7
+ ua = -3.572492586e-09 lua = 2.469456457e-16 wua = 1.978629571e-14 pua = -3.922422012e-21
+ ub = 4.262535660e-18 lub = -1.687925808e-25 wub = -1.950403152e-23 pub = 3.184917676e-30
+ uc = -2.180019591e-11 luc = 1.473801867e-17 wuc = 7.669034579e-16 puc = -1.647843525e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.178462721e-03 lu0 = 4.698216784e-09 wu0 = 1.844666042e-07 pu0 = -4.203558945e-14
+ a0 = 7.577763427e+00 la0 = -1.444321709e-06 wa0 = -1.082144394e-05 pa0 = 2.062567215e-12
+ keta = 8.184019325e-01 lketa = -1.942150896e-07 wketa = -3.553778092e-06 pketa = 7.865837251e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.359754981e+00 lags = 8.755521481e-07 wags = 5.643185463e-07 pags = -1.470614132e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.899302647e-01 lvoff = 2.230304255e-08 wvoff = 9.597306212e-08 pvoff = -3.465739477e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.333966648e+00 lnfactor = 3.227810349e-07 wnfactor = 5.374355517e-06 pnfactor = -9.584523694e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.302623816e-06 lcit = 1.642463767e-12 wcit = 4.338505643e-11 pcit = -1.130614571e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -7.560291898e-02 leta0 = 2.264813803e-08 weta0 = -7.831815720e-07 peta0 = 1.941720327e-13
+ etab = 1.964671272e-01 letab = -3.922923143e-08 wetab = -1.774131531e-06 petab = 3.309664682e-13
+ dsub = -5.509021671e-01 ldsub = 1.682484483e-07 wdsub = 4.681982856e-06 pdsub = -9.054050933e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.185564234e-01 lpclm = -1.223875514e-07 wpclm = 1.326954952e-06 ppclm = -2.897974907e-13
+ pdiblc1 = -1.270952915e+00 lpdiblc1 = 4.328443297e-07 wpdiblc1 = 6.923572081e-11 ppdiblc1 = -1.804282884e-17
+ pdiblc2 = -1.920896613e-02 lpdiblc2 = 7.996026579e-09 wpdiblc2 = 2.325599289e-07 ppdiblc2 = -5.617993145e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.423466313e-02 lalpha0 = -4.897488775e-09 walpha0 = -1.055168547e-07 palpha0 = 2.287204265e-14
+ alpha1 = 0.0
+ beta0 = 5.429419371e+01 lbeta0 = -5.491968223e-06 wbeta0 = -1.159664388e-04 pbeta0 = 2.672008248e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.865147651e-01 lkt1 = 1.169363632e-08 wkt1 = 1.545276520e-06 pkt1 = -2.792931040e-13
+ kt2 = -1.051028938e-01 lkt2 = 2.458256332e-08 wkt2 = 4.612179405e-07 pkt2 = -1.396959844e-13
+ at = 7.102537653e+04 lat = 2.040153817e-04 wat = -5.722142389e-01 pat = 1.193545486e-7
+ ute = -6.648105127e+00 lute = 7.523422088e-07 wute = 3.872588465e-05 pute = -6.335504544e-12
+ ua1 = -1.564436843e-08 lua1 = 2.855163019e-15 wua1 = 1.199111170e-13 pua1 = -2.195925965e-20
+ ub1 = 1.306814430e-17 lub1 = -2.490413500e-24 wub1 = -1.056748562e-22 pub1 = 1.998033207e-29
+ uc1 = -4.982853807e-10 luc1 = 9.624047388e-17 wuc1 = 2.458365668e-15 puc1 = -4.748168139e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.15 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.468756752e-01 lvth0 = 6.820892244e-08 wvth0 = 1.788186980e-06 pvth0 = -2.728536138e-13
+ k1 = 1.828459196e+00 lk1 = -2.178257973e-07 wk1 = -5.033482715e-06 pk1 = 9.763113620e-13
+ k2 = -3.804817216e-01 lk2 = 5.303830422e-08 wk2 = 1.199837101e-06 pk2 = -2.528749141e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.382701899e+05 lvsat = -2.477426968e-02 wvsat = -7.611935348e-01 pvsat = 1.268991525e-7
+ ua = -7.860820927e-09 lua = 1.064301028e-15 wua = 2.800053283e-14 pua = -5.488055609e-21
+ ub = 1.628561958e-17 lub = -2.460392375e-24 wub = -7.115549826e-23 pub = 1.302968724e-29
+ uc = 5.039079882e-10 luc = -8.546196121e-17 wuc = -1.911166624e-15 puc = 3.456558051e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.632265940e-02 lu0 = -6.261497093e-09 wu0 = -2.363129607e-07 pu0 = 3.816499562e-14
+ a0 = 0.0
+ keta = 8.080350157e-01 lketa = -1.922391553e-07 wketa = -3.962649485e-06 pketa = 8.645146125e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.151353997e+00 lags = 1.573477678e-08 wags = -1.382007447e-06 pags = 2.239083211e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -5.093335580e-01 lvoff = 8.318131024e-08 wvoff = 2.620210109e-06 pvoff = -5.157769759e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -4.017490158e+00 lnfactor = 1.342768702e-06 wnfactor = 2.612273825e-05 pnfactor = -4.913094119e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.970612224e-05 lcit = -2.361803231e-12 wcit = -1.012317983e-10 pcit = 1.625782681e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -4.024696278e-01 leta0 = 8.494893274e-08 weta0 = 3.217482977e-06 peta0 = -5.683546303e-13
+ etab = -2.198226399e-01 letab = 4.011559818e-08 wetab = 8.647229346e-07 petab = -1.719991930e-13
+ dsub = 7.163498423e-01 ldsub = -7.328978467e-08 wdsub = -4.339720272e-07 pdsub = 6.969590756e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.677148020e+00 lpclm = -2.860351097e-07 wpclm = -1.106370759e-05 ppclm = 2.071862790e-12
+ pdiblc1 = 1.110385018e+01 lpdiblc1 = -1.925793140e-06 wpdiblc1 = -4.687328981e-05 ppdiblc1 = 8.934044192e-12
+ pdiblc2 = 1.548168627e-01 lpdiblc2 = -2.517329639e-08 wpdiblc2 = -5.234523186e-07 ppdiblc2 = 8.791600293e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.984633136e-03 lalpha0 = 1.243509092e-09 walpha0 = 6.855570983e-08 palpha0 = -1.030618815e-14
+ alpha1 = 0.0
+ beta0 = 1.903818858e+01 lbeta0 = 1.227826354e-06 wbeta0 = 8.824422678e-05 pbeta0 = -1.220247038e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 2.000206238e-01 lkt1 = -1.001000088e-07 wkt1 = -3.373466848e-06 pkt1 = 6.582193820e-13
+ kt2 = 4.504385310e-01 lkt2 = -8.130363225e-08 wkt2 = -2.884793785e-06 pkt2 = 4.980538504e-13
+ at = -1.158710764e+05 lat = 3.582647931e-02 wat = 1.207487730e+00 pat = -2.198566467e-7
+ ute = -4.688617754e+00 lute = 3.788639155e-07 wute = 1.094031175e-05 pute = -1.039574348e-12
+ ua1 = -8.508617133e-09 lua1 = 1.495088821e-15 wua1 = 3.721524752e-14 pua1 = -6.197426918e-21
+ ub1 = 7.554705620e-18 lub1 = -1.439552088e-24 wub1 = -3.031955146e-23 pub1 = 5.617610989e-30
+ uc1 = -3.280166061e-10 luc1 = 6.378724544e-17 wuc1 = 2.300157716e-15 puc1 = -4.446623781e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.16 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.431261
+ k1 = 0.40031
+ k2 = -0.007143591
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 242950.0
+ ua = -1.26631373e-9
+ ub = 2.614475e-18
+ uc = 7.0441e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03251371
+ a0 = 1.928858
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.527887
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11890341
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.05278474
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.068446
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25403
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.17 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.431261
+ k1 = 0.40031
+ k2 = -0.007143591
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 242950.0
+ ua = -1.26631373e-9
+ ub = 2.614475e-18
+ uc = 7.0441e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03251371
+ a0 = 1.928858
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.527887
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11890341
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.05278474
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.068446
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25403
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.18 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.375025056e-01 lvth0 = -2.503218228e-8
+ k1 = 3.048266060e-01 lk1 = 3.829457000e-7
+ k2 = 2.784367289e-02 lk2 = -1.403199205e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.383139702e+05 lvsat = -7.835267389e-1
+ ua = -1.280239276e-09 lua = 5.584979595e-17
+ ub = 2.675408244e-18 lub = -2.443788668e-25
+ uc = 4.442584660e-11 luc = 1.043363742e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.216794712e-02 lu0 = 1.386716615e-9
+ a0 = 1.947956689e+00 la0 = -7.659720371e-8
+ keta = 2.171448000e-01 lketa = -8.708809349e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.177341639e-01 lags = 3.391448240e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.264962398e-01 lvoff = 3.045180336e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.345022689e-01 lnfactor = 2.479683679e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.502650000e-05 lcit = -2.015928090e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 6.993782904e-01 ldsub = -5.589905717e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.768744200e-02 lpclm = -7.716972729e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.378959080e-03 lpdiblc2 = 8.855568914e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.202347795e-05 lalpha0 = 3.842693261e-10 palpha0 = 1.262177448e-29
+ alpha1 = 0.0
+ beta0 = 1.374529394e+01 lbeta0 = 1.522448650e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.434039790e-01 lkt1 = -4.261671982e-8
+ kt2 = -4.760006260e-02 lkt2 = 5.177709706e-8
+ at = 7.801228450e+04 lat = -3.977426122e-2
+ ute = -1.160206550e+00 lute = -1.471627506e-7
+ ua1 = 3.222567210e-09 lua1 = -1.192219872e-15
+ ub1 = -3.672807280e-18 lub1 = 1.603066017e-24
+ uc1 = -1.439063870e-11 luc1 = -5.048287123e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.19 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.138036135e-01 lvth0 = 2.261681010e-8
+ k1 = 5.556228200e-01 lk1 = -1.213051679e-07 wk1 = -5.421010862e-20
+ k2 = -5.979197904e-02 lk2 = 3.588032122e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.297101440e+04 lvsat = 5.156180805e-2
+ ua = -9.689957784e-10 lua = -5.699363808e-16
+ ub = 2.444872822e-18 lub = 2.191356523e-25
+ uc = 1.166795582e-10 luc = -4.093693832e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.615508621e-02 lu0 = -6.629825244e-9
+ a0 = 2.062631391e+00 la0 = -3.071621595e-7
+ keta = -2.633870340e-01 lketa = 9.527637056e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.254696020e-01 lags = 1.293982748e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.071038869e-01 lvoff = -8.538461481e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.575622568e+00 lnfactor = 1.853472052e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.277005460e-04 leta0 = -5.569471779e-11
+ etab = -5.239310080e-04 letab = 4.811568468e-11
+ dsub = -1.634205809e-01 ldsub = 1.175752839e-06 pdsub = -5.169878828e-26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.771532904e-01 lpclm = 4.553190493e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.505417840e-03 lpdiblc2 = 6.590710931e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.991262076e-04 lalpha0 = -1.407982317e-10
+ alpha1 = 0.0
+ beta0 = 2.140035606e+01 lbeta0 = -1.667813984e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.647819080e-01 lkt1 = 3.657442248e-10
+ kt2 = -7.919910800e-03 lkt2 = -2.800381615e-8
+ at = 4.254043500e+04 lat = 3.154543939e-2
+ ute = -1.294642360e+00 lute = 1.231338890e-7
+ ua1 = 3.087603920e-09 lua1 = -9.208626816e-16
+ ub1 = -3.599190660e-18 lub1 = 1.455052441e-24 wub1 = 3.761581923e-37
+ uc1 = -5.101882940e-11 luc1 = 2.316176899e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.20 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.426783384e-01 lvth0 = -6.563986827e-9
+ k1 = 4.270119200e-01 lk1 = 8.669007648e-9
+ k2 = -1.654236752e-02 lk2 = -7.827736185e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -5.747626680e+04 lvsat = 1.328618304e-01 pvsat = -6.776263578e-21
+ ua = -1.441970692e-09 lua = -9.194793282e-17
+ ub = 2.774930444e-18 lub = -1.144205807e-25
+ uc = 9.694299559e-11 luc = -2.099116814e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.120788752e-02 lu0 = -1.630186248e-9
+ a0 = 1.956386129e+00 la0 = -1.997906976e-7
+ keta = -3.418051320e-01 lketa = 1.745257004e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.001181235e+00 lags = -2.016451428e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.166392140e-01 lvoff = 1.097940139e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.423125243e+00 lnfactor = 3.394610015e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.551990035e-04 leta0 = -4.877245624e-10
+ etab = -8.983088033e-04 letab = 4.264618846e-10
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.597508640e-01 lpclm = 1.148437108e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.421073408e-02 lpdiblc2 = -2.206881661e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.299440988e-06 lalpha0 = 6.175192876e-11
+ alpha1 = 0.0
+ beta0 = 1.847349677e+01 lbeta0 = 2.791102599e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.632558320e-01 lkt1 = -1.176508181e-9
+ kt2 = -3.686054600e-02 lkt2 = 1.243589788e-9
+ at = 9.774298800e+04 lat = -2.424226067e-2
+ ute = -1.303717840e+00 lute = 1.323055691e-7
+ ua1 = 1.943566400e-09 lua1 = 2.353016362e-16
+ ub1 = -1.756332360e-18 lub1 = -4.073401570e-25
+ uc1 = -3.018733280e-11 luc1 = 2.109458528e-18 wuc1 = 3.155443621e-30
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.21 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.600650913e-02 lvth0 = 2.378524963e-07 wvth0 = 2.616917201e-06 pvth0 = -1.336197923e-12
+ k1 = 2.800830240e-01 lk1 = 8.369090195e-8
+ k2 = 6.497932819e-02 lk2 = -4.945271402e-08 wk2 = -1.944114756e-07 pk2 = 9.926649944e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.356249646e+04 lvsat = 1.155454593e-01 wvsat = 1.236702718e+00 pvsat = -6.314604078e-7
+ ua = -1.134656613e-08 lua = 4.965338495e-15 wua = 4.819925776e-14 pua = -2.461054101e-20
+ ub = 1.144221286e-17 lub = -4.539934984e-24 wub = -4.174750727e-23 pub = 2.131627721e-29
+ uc = 4.937028284e-11 luc = 3.299458988e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -6.081337997e-02 lu0 = 4.535587293e-08 wu0 = 4.715243060e-07 pu0 = -2.407603106e-13
+ a0 = 1.688937120e+00 la0 = -6.323123347e-8
+ keta = 3.688404081e-02 lketa = -1.883299124e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.062068424e-01 lags = -2.767750313e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.172397928e-01 lvoff = 1.404595627e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.175698395e+01 lnfactor = 7.069224757e-06 wnfactor = 6.404532759e-05 pnfactor = -3.270154427e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -3.737219299e-03 leta0 = 1.908224365e-9
+ etab = 5.850190428e-02 letab = -2.990328692e-08 wetab = 1.111730743e-21 petab = -3.534096855e-28
+ dsub = 1.688504919e+00 ldsub = -3.515506114e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.765288560e-01 lpclm = 4.156868126e-9
+ pdiblc1 = 0.39
+ pdiblc2 = 4.648038240e-03 lpdiblc2 = 2.675830835e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.677617963e-03 lalpha0 = 9.176801660e-10 walpha0 = -2.646977960e-23 palpha0 = -2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.710456674e+01 lbeta0 = 3.490078270e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.863037600e-01 lkt1 = 1.059176386e-8
+ kt2 = -4.326872160e-02 lkt2 = 4.515604249e-9
+ at = 5.194013680e+04 lat = -8.553248501e-4
+ ute = -1.258458784e+00 lute = 1.091962951e-7
+ ua1 = 2.266177760e-09 lua1 = 7.057627574e-17
+ ub1 = -2.748924560e-18 lub1 = 9.947742034e-26
+ uc1 = -5.321677440e-11 luc1 = 1.386829141e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.22 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 2.492528357e+00 lvth0 = -4.210836899e-07 wvth0 = -9.346132862e-06 pvth0 = 1.781372923e-12
+ k1 = 3.224366571e-01 lk1 = 7.265354515e-8
+ k2 = -1.162191978e-01 lk2 = -2.232378139e-09 wk2 = 6.943266986e-07 pk2 = -1.323386687e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.048440307e+06 lvsat = -1.638184714e-01 wvsat = -4.416795421e+00 pvsat = 8.418412073e-7
+ ua = 3.532903103e-08 lua = -7.198322123e-15 wua = -1.721402063e-13 pua = 3.280992332e-20
+ ub = -2.991140691e-17 lub = 6.236818329e-24 wub = 1.490982402e-22 pub = -2.841812459e-29
+ uc = 1.336432299e-10 luc = -1.866207102e-17 wuc = 1.262177448e-29
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.775435753e-01 lu0 = -6.887994960e-08 wu0 = -1.684015379e-06 pu0 = 3.209733311e-13
+ a0 = 5.384368286e+00 la0 = -1.026260595e-6
+ keta = 9.808774473e-02 lketa = -3.478267648e-08 pketa = 1.615587134e-27
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.245373429e+00 lags = 8.457443155e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.704775143e-01 lvoff = 1.527834587e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.878517789e+01 lnfactor = -8.708062620e-06 wnfactor = -2.287333128e-04 pnfactor = 4.359656943e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 7.491079919e-06 lcit = -6.491754269e-13
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.343457508e-01 leta0 = 6.200480756e-08 peta0 = 1.615587134e-27
+ etab = -1.631310468e-01 letab = 2.785426014e-08 wetab = -1.355252716e-20
+ dsub = 3.980874970e-01 ldsub = -1.526783136e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.087516514e+00 lpclm = -1.811265156e-7
+ pdiblc1 = -1.270938882e+00 lpdiblc1 = 4.328406726e-7
+ pdiblc2 = 2.792853429e-02 lpdiblc2 = -3.391066435e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.847484325e-03 lalpha0 = -2.615614903e-10
+ alpha1 = 0.0
+ beta0 = 3.078899191e+01 lbeta0 = -7.608292872e-8
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -7.330314286e-02 lkt1 = -4.491619697e-8
+ kt2 = -1.161877143e-02 lkt2 = -3.732372766e-9
+ at = -4.495655143e+04 lat = 2.439595210e-2
+ ute = 1.201232514e+00 lute = -5.317992572e-7
+ ua1 = 8.660378971e-09 lua1 = -1.595752560e-15
+ ub1 = -8.351059771e-18 lub1 = 1.559393856e-24
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.23 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -7.386775378e-01 lvth0 = 1.947841537e-07 wvth0 = 4.707930239e-06 pvth0 = -8.973315036e-13
+ k1 = 8.082241333e-01 lk1 = -1.993754781e-8
+ k2 = -4.102284470e-01 lk2 = 5.380578475e-08 wk2 = 1.346597033e-06 pk2 = -2.566613945e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.385330472e+04 lvsat = 2.765581132e-02 wvsat = 6.913563310e-01 pvsat = -1.317725167e-7
+ ua = -1.301021841e-08 lua = 2.015138821e-15 wua = 5.340585774e-14 pua = -1.017915649e-20
+ ub = -1.420528542e-18 lub = 8.064569121e-25 wub = 1.620043940e-23 pub = -3.087803749e-30
+ uc = 1.165342133e-10 luc = -1.540109246e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -9.635991765e-02 lu0 = 2.144605615e-08 wu0 = 5.169694356e-07 pu0 = -9.853437442e-14
+ a0 = 0.0
+ keta = 4.846811240e-03 lketa = -1.701095456e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 8.712353333e-01 lags = 6.111868547e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = 2.175602256e-02 lvoff = -2.136136626e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -8.269658632e+01 lnfactor = 1.635236164e-05 wnfactor = 4.142978611e-04 pnfactor = -7.896517232e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -8.125198107e-07 lcit = 9.334906816e-13
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.496810064e-01 leta0 = -3.025069235e-8
+ etab = -4.455221445e-02 letab = 5.253134690e-9
+ dsub = 6.283881857e-01 ldsub = -5.916314262e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.653514667e-01 lpclm = 1.339101215e-7
+ pdiblc1 = 1.603117493e+00 lpdiblc1 = -1.149544725e-7
+ pdiblc2 = 4.871847333e-02 lpdiblc2 = -7.353628817e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.910902588e-03 lalpha0 = -8.454490111e-10
+ alpha1 = 0.0
+ beta0 = 3.692438375e+01 lbeta0 = -1.245488613e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.837463333e-01 lkt1 = 3.331427513e-8
+ kt2 = -1.342794333e-01 lkt2 = 1.964674939e-08 wkt2 = -1.355252716e-20
+ at = 1.288742400e+05 lat = -8.736196744e-3
+ ute = -2.471129333e+00 lute = 1.681529109e-7
+ ua1 = -9.654700667e-10 lua1 = 2.389342667e-16
+ ub1 = 1.409245067e-18 lub1 = -3.009202457e-25 pub1 = 1.121038771e-44
+ uc1 = 1.382016533e-10 luc1 = -2.634123513e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.24 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.396315006e-01 wvth0 = -4.087859533e-8
+ k1 = 2.494330533e-01 wk1 = 7.368302009e-7
+ k2 = 5.272278487e-02 wk2 = -2.923664265e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.493316251e+05 wvsat = -5.195306235e-1
+ ua = -1.506061110e-09 wua = 1.170842292e-15
+ ub = 2.915846466e-18 wub = -1.471792762e-24
+ uc = 7.252139330e-11 wuc = -1.015991275e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.257610524e-02 wu0 = -3.047164989e-10
+ a0 = 2.284318619e+00 wa0 = -1.735945252e-6
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.124209497e-01 wags = 7.553077663e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.248638928e-01 wvoff = 2.910891169e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 5.307523946e-01 wnfactor = 2.549423263e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.727047739e-05 wcit = -3.550646689e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.228460764e-01 wpclm = 9.342035491e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 6.405965113e-03 wpdiblc2 = 8.841110256e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.647008226e-05 walpha0 = 3.574766232e-11
+ alpha1 = 0.0
+ beta0 = 1.717144284e+01 wbeta0 = 1.806526428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.514562510e-01 wkt1 = -1.256928928e-8
+ kt2 = -3.455913141e-02 wkt2 = -6.391164040e-10
+ at = -2.959886961e+05 wat = 1.778057342e+0
+ ute = -1.103692480e+00 wute = -4.551929055e-7
+ ua1 = 4.147321839e-09 wua1 = -5.967926955e-15
+ ub1 = -4.995330683e-18 wub1 = 8.410771877e-24
+ uc1 = 1.877070653e-12 wuc1 = -1.409180658e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.25 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.396315006e-01 wvth0 = -4.087859533e-8
+ k1 = 2.494330533e-01 wk1 = 7.368302009e-7
+ k2 = 5.272278487e-02 wk2 = -2.923664265e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.493316251e+05 wvsat = -5.195306235e-1
+ ua = -1.506061110e-09 wua = 1.170842292e-15
+ ub = 2.915846466e-18 wub = -1.471792762e-24
+ uc = 7.252139330e-11 wuc = -1.015991275e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.257610524e-02 wu0 = -3.047164989e-10
+ a0 = 2.284318619e+00 wa0 = -1.735945252e-6
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.124209497e-01 wags = 7.553077663e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.248638928e-01 wvoff = 2.910891169e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 5.307523946e-01 wnfactor = 2.549423263e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.727047739e-05 wcit = -3.550646689e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.228460764e-01 wpclm = 9.342035491e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 6.405965113e-03 wpdiblc2 = 8.841110256e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.647008226e-05 walpha0 = 3.574766232e-11
+ alpha1 = 0.0
+ beta0 = 1.717144284e+01 wbeta0 = 1.806526428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.514562510e-01 wkt1 = -1.256928928e-8
+ kt2 = -3.455913141e-02 wkt2 = -6.391164040e-10
+ at = -2.959886961e+05 wat = 1.778057342e+0
+ ute = -1.103692480e+00 wute = -4.551929055e-7
+ ua1 = 4.147321839e-09 wua1 = -5.967926955e-15
+ ub1 = -4.995330683e-18 wub1 = 8.410771877e-24
+ uc1 = 1.877070653e-12 wuc1 = -1.409180658e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.26 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.688440581e-01 lvth0 = -1.171598829e-07 wvth0 = -1.530611728e-07 pvth0 = 4.499194452e-13
+ k1 = -7.492470859e-02 lk1 = 1.300869240e-06 wk1 = 1.854572508e-06 pk1 = -4.482817295e-12
+ k2 = 1.820446314e-01 lk2 = -5.186581976e-07 wk2 = -7.530635110e-07 pk2 = 1.847671727e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.362877347e+05 lvsat = -1.150866173e+00 wvsat = -9.668345752e-01 pvsat = 1.793957228e-6
+ ua = -1.736282479e-09 lua = 9.233258244e-16 wua = 2.227155389e-15 pua = -4.236449307e-21
+ ub = 3.277098198e-18 lub = -1.448836194e-24 wub = -2.938443144e-24 pub = 5.882148025e-30
+ uc = 3.777155232e-11 luc = 1.393677122e-16 wuc = 3.249724426e-17 puc = -1.710807939e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.149368176e-02 lu0 = 4.341167586e-09 wu0 = 3.292876003e-09 pu0 = -1.442850449e-14
+ a0 = 2.531747594e+00 la0 = -9.923386451e-07 wa0 = -2.851030449e-06 pa0 = 4.472160690e-12
+ keta = 1.647976638e-01 lketa = -6.609375105e-07 wketa = 2.556450916e-07 pketa = -1.025290205e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.976295675e-01 lags = 1.262502317e-06 wags = -2.516856087e-06 pags = 1.039702675e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.480268893e-01 lvoff = 9.289751387e-08 wvoff = 1.051481562e-07 pvoff = -3.049629941e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.113825429e+00 lnfactor = 6.595743820e-06 wnfactor = 7.561490562e-06 pnfactor = -2.010139711e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.960598830e-05 lcit = -4.947280008e-11 wcit = -7.120111806e-11 pcit = 1.431569680e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398569041e-01 letab = 2.801680995e-07 wetab = -5.589782372e-11 petab = 2.241838118e-16
+ dsub = 5.866338881e-01 ldsub = -1.068178715e-07 wdsub = 5.506042007e-07 pdsub = -2.208253207e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -9.936540810e-02 lpclm = -9.417156841e-08 wpclm = 9.135006514e-07 ppclm = 8.303104142e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 2.846049534e-03 lpdiblc2 = 1.427739742e-08 wpdiblc2 = 7.486193705e-09 ppdiblc2 = -2.647831279e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.782516840e-05 lalpha0 = 3.380745323e-10 walpha0 = -2.050307442e-11 palpha0 = 2.255992048e-16
+ alpha1 = 0.0
+ beta0 = 1.322558698e+01 lbeta0 = 1.582524948e-05 wbeta0 = 2.538066886e-06 pbeta0 = -2.933916164e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.219583638e-01 lkt1 = -1.183042264e-07 wkt1 = -1.047328786e-07 pkt1 = 3.696312913e-13
+ kt2 = -6.838465965e-02 lkt2 = 1.356606636e-07 wkt2 = 1.015046974e-07 pkt2 = -4.096579795e-13
+ at = -6.747470705e+05 lat = 1.519048337e+00 wat = 3.676213224e+00 pat = -7.612743980e-6
+ ute = -9.395298795e-01 lute = -6.583905251e-07 wute = -1.077707622e-06 pute = 2.496657521e-12
+ ua1 = 5.086904929e-09 lua1 = -3.768291938e-15 wua1 = -9.104772899e-15 pua1 = 1.258063434e-20
+ ub1 = -6.577051209e-18 lub1 = 6.343648340e-24 wub1 = 1.418331086e-23 pub1 = -2.315134486e-29
+ uc1 = 2.302620734e-11 luc1 = -8.482072760e-17 wuc1 = -1.827307802e-16 puc1 = 1.676940723e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.27 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.863920332e-01 lvth0 = 4.861815826e-08 wvth0 = 1.338685642e-07 pvth0 = -1.269814840e-13
+ k1 = 7.131484205e-01 lk1 = -2.836305937e-07 wk1 = -7.692998991e-07 pk1 = 7.927405659e-13
+ k2 = -1.265747776e-01 lk2 = 1.018519861e-07 wk2 = 3.261438144e-07 pk2 = -3.221825214e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.978344050e+04 lvsat = 8.253360795e-03 wvsat = -1.797790047e-01 pvsat = 2.115032984e-7
+ ua = -9.537569882e-10 lua = -6.500199281e-16 wua = -7.442091797e-17 pua = 3.911000156e-22
+ ub = 2.214939918e-18 lub = 6.867392441e-25 wub = 1.122911827e-24 pub = -2.283612281e-30
+ uc = 1.344390431e-10 luc = -5.499194470e-17 wuc = -8.673110840e-17 puc = 6.863973193e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.512322968e-02 lu0 = -2.956401448e-09 wu0 = 5.039226164e-09 pu0 = -1.793971612e-14
+ a0 = 1.995617801e+00 la0 = 8.560391543e-08 wa0 = 3.272709196e-07 pa0 = -1.918132042e-12
+ keta = -1.827045369e-01 lketa = 3.775041422e-08 wketa = -3.940250771e-07 pketa = 2.809366367e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.976885917e-01 lags = 2.258389008e-06 wags = 4.996746513e-06 pags = -4.709822632e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -8.875202117e-02 lvoff = -2.628053598e-08 wvoff = -8.962408901e-08 pvoff = 8.664608212e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.807009285e+00 lnfactor = -1.287486457e-06 wnfactor = -6.013661742e-06 pnfactor = 7.192804115e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.177372757e-04 leta0 = -3.566256658e-11 weta0 = 4.865712486e-11 peta0 = -9.783001524e-17
+ etab = -5.415766835e-04 letab = 6.070225757e-11 wetab = 8.617530295e-11 petab = -6.146841665e-17
+ dsub = -2.534808307e-01 ldsub = 1.582316782e-06 wdsub = 4.398227389e-07 pdsub = -1.985516000e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.396780468e-01 lpclm = 1.394301023e-06 wpclm = 3.235539027e-06 ppclm = -4.585659316e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 9.610058591e-03 lpdiblc2 = 6.776808117e-10 wpdiblc2 = -2.004562880e-08 ppdiblc2 = 2.887716954e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.429512492e-04 lalpha0 = -6.560653286e-11 walpha0 = 2.743388360e-10 palpha0 = -3.672099403e-16
+ alpha1 = 0.0
+ beta0 = 2.033465129e+01 lbeta0 = 1.531764794e-06 wbeta0 = 5.204529110e-06 pbeta0 = -8.295105110e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.984823825e-01 lkt1 = 3.555496559e-08 wkt1 = 1.645813222e-07 pkt1 = -1.718518409e-13
+ kt2 = 5.574947439e-02 lkt2 = -1.139234263e-07 wkt2 = -3.109389930e-07 pkt2 = 4.196013043e-13
+ at = 9.282907453e+04 lat = -2.424026075e-02 wat = -2.455921144e-01 pat = 2.724378345e-7
+ ute = -1.264455280e+00 lute = -5.095515458e-09 wute = -1.474231346e-07 pute = 6.262275312e-13
+ ua1 = 5.028816322e-09 lua1 = -3.651498986e-15 wua1 = -9.480201947e-15 pua1 = 1.333547199e-20
+ ub1 = -6.020880034e-18 lub1 = 5.225410576e-24 wub1 = 1.182668331e-23 pub1 = -1.841310950e-29
+ uc1 = -9.789132403e-11 luc1 = 1.582960610e-16 wuc1 = 2.289088584e-16 puc1 = -6.599485851e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.28 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.462953823e-01 lvth0 = -1.192016635e-08 wvth0 = -1.766437675e-08 pvth0 = 2.615770613e-14
+ k1 = 4.013290284e-01 lk1 = 3.149408394e-08 wk1 = 1.254262534e-07 pk1 = -1.114696838e-13
+ k2 = -1.454307333e-02 lk2 = -1.136725423e-08 wk2 = -9.763853059e-09 pk2 = 1.728576730e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -9.163355237e+04 lvsat = 1.612753738e-01 wvsat = 1.668122277e-01 pvsat = -1.387618010e-7
+ ua = -1.034320785e-09 lua = -5.686021551e-16 wua = -1.990819471e-15 pua = 2.327812393e-21
+ ub = 2.583603010e-18 lub = 3.141683229e-25 wub = 9.343762224e-25 pub = -2.093078199e-30
+ uc = 9.363132046e-11 luc = -1.375166021e-17 wuc = 1.617306223e-17 puc = -3.535522291e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.813730840e-02 lu0 = -6.002429405e-09 wu0 = -3.384086627e-08 pu0 = 2.135250529e-14
+ a0 = 2.964782162e+00 la0 = -8.938335876e-07 wa0 = -4.924653286e-06 pa0 = 3.389462560e-12
+ keta = -3.117534833e-01 lketa = 1.681672794e-07 wketa = -1.467617344e-07 pketa = 3.105230257e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.984823776e+00 lags = -3.080117991e-06 wags = -4.803765898e-06 pags = 5.194575210e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.100549538e-01 lvoff = -4.751792266e-09 wvoff = -3.215522253e-08 pvoff = 2.856804566e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.562156034e+00 lnfactor = -2.943776145e-08 wnfactor = -6.789777215e-07 pnfactor = 1.801572444e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.899747706e-04 leta0 = -5.129056788e-10 weta0 = -1.698326577e-10 peta0 = 1.229757590e-16
+ etab = -9.627047148e-04 letab = 4.862942460e-10 wetab = 3.144870931e-10 petab = -2.922003118e-16
+ dsub = 1.631098109e+00 ldsub = -3.222386945e-07 wdsub = -3.082062281e-06 pdsub = 1.573701000e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.642046070e-01 lpclm = -2.446278698e-08 wpclm = -1.975210522e-06 ppclm = 6.803241781e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.220658290e-02 lpdiblc2 = -1.946366655e-09 wpdiblc2 = 9.787572910e-09 ppdiblc2 = -1.272264110e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.070122836e-05 lalpha0 = 5.793933817e-11 walpha0 = -1.074435689e-10 palpha0 = 1.861935806e-17
+ alpha1 = 0.0
+ beta0 = 1.942818654e+01 lbeta0 = 2.447838063e-06 wbeta0 = -4.662370716e-06 pbeta0 = 1.676383854e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.503310462e-01 lkt1 = -1.310677488e-08 wkt1 = -6.312013024e-08 pkt1 = 5.826324697e-14
+ kt2 = -6.589998840e-02 lkt2 = 9.015520761e-09 wkt2 = 1.418184729e-07 pkt2 = -3.795539070e-14
+ at = 1.198833680e+05 lat = -5.158132970e-02 wat = -1.081258666e-01 pat = 1.335144444e-7
+ ute = -2.238208352e+00 lute = 9.789793391e-07 wute = 4.563724588e-06 pute = -4.134858357e-12
+ ua1 = -2.726467352e-09 lua1 = 4.185990695e-15 wua1 = 2.280681033e-14 pua1 = -1.929378262e-20
+ ub1 = 4.584300525e-18 lub1 = -5.492184897e-24 wub1 = -3.096543179e-23 pub1 = 2.483260202e-29
+ uc1 = 1.840337005e-10 luc1 = -1.266173688e-16 wuc1 = -1.046180549e-15 puc1 = 6.286567704e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.29 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.986357867e-01 lvth0 = -3.864517681e-08 wvth0 = 5.911353450e-09 pvth0 = 1.411993829e-14
+ k1 = 3.022304018e-01 lk1 = 8.209384270e-08 wk1 = -1.081600416e-07 pk1 = 7.799478407e-15
+ k2 = 2.269182158e-02 lk2 = -3.037939157e-08 wk2 = 1.210590608e-08 pk2 = 6.119068285e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.831693614e+05 lvsat = -3.009899396e-02 wvsat = -2.612683195e-01 pvsat = 7.981612636e-8
+ ua = -3.334837986e-09 lua = 6.060419277e-16 wua = 9.072781630e-15 pua = -3.321262329e-21
+ ub = 4.771594755e-18 lub = -8.030202619e-25 wub = -9.170543144e-24 pub = 3.066493629e-30
+ uc = 4.954613784e-11 luc = 8.758234036e-18 wuc = -8.588142757e-19 puc = -2.665874676e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.453324036e-02 lu0 = 9.438077358e-10 wu0 = 5.472128360e-08 pu0 = -2.386732843e-14
+ a0 = 1.045429869e+00 la0 = 8.618769327e-08 wa0 = 3.142664187e-06 pa0 = -7.297097416e-13
+ keta = 7.608545142e-02 lketa = -2.986328062e-08 wketa = -1.914459690e-07 pketa = 5.386807273e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.139467883e+00 lags = 5.575453303e-07 wags = 1.096708937e-05 pags = -2.858023490e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.254556026e-01 lvoff = 3.111779014e-09 wvoff = 4.012313980e-08 pvoff = -8.337286147e-15
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -2.786158941e-01 lnfactor = 9.104603851e-07 wnfactor = 7.988995421e-06 pnfactor = -2.624294643e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.238031453e-03 leta0 = -1.660763306e-09 weta0 = -3.406468358e-08 peta0 = 1.742968664e-14
+ etab = 1.156574142e-01 letab = -5.905993846e-08 wetab = -2.791275059e-07 petab = 1.423908813e-13
+ dsub = 1.574327190e+00 ldsub = -2.932514631e-07 wdsub = 5.576040647e-07 pdsub = -2.847126354e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.996401639e-01 lpclm = -4.255618234e-08 wpclm = -1.089597539e-06 ppclm = 2.281301889e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 4.902668738e-03 lpdiblc2 = 1.783011916e-09 wpdiblc2 = -1.243526231e-09 ppdiblc2 = 4.360215111e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.396392408e-03 lalpha0 = 7.815073487e-10 walpha0 = -1.373407182e-09 palpha0 = 6.650203792e-16
+ alpha1 = 0.0
+ beta0 = 1.764033415e+01 lbeta0 = 3.360715495e-06 wbeta0 = -2.616500484e-06 pbeta0 = 6.317625134e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.460514846e-01 lkt1 = 3.576808097e-08 wkt1 = 2.917869752e-07 pkt1 = -1.229523211e-13
+ kt2 = -6.032463105e-02 lkt2 = 6.168743301e-09 wkt2 = 8.329509220e-08 pkt2 = -8.073352529e-15
+ at = -4.768550074e+02 lat = 9.874600155e-03 wat = 2.559862420e-01 pat = -5.240119825e-8
+ ute = -1.072179475e+00 lute = 3.836049946e-07 wute = -9.097229479e-07 pute = -1.340116045e-12
+ ua1 = 4.705219949e-09 lua1 = 3.913711593e-16 wua1 = -1.191142839e-14 pua1 = -1.566649933e-21
+ ub1 = -6.455251943e-18 lub1 = 1.446105931e-25 wub1 = 1.810040573e-23 pub1 = -2.204146190e-31
+ uc1 = -1.763003973e-10 luc1 = 5.736922150e-17 wuc1 = 6.010973348e-16 puc1 = -2.124433172e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.30 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 6.226325442e-01 lvth0 = -7.095873181e-08 wvth0 = -2.142161733e-07 pvth0 = 7.148517175e-14
+ k1 = 3.376497671e-01 lk1 = 7.286355611e-08 wk1 = -7.429550421e-08 pk1 = -1.025620028e-15
+ k2 = 1.583106600e-02 lk2 = -2.859147867e-08 wk2 = 4.943942772e-08 pk2 = -3.610047456e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.902217631e+04 lvsat = 1.788976246e-02 wvsat = 2.198304345e-01 pvsat = -4.555820893e-8
+ ua = 3.581993886e-09 lua = -1.196484458e-15 wua = -1.709878833e-14 pua = 3.499048803e-21
+ ub = -2.255406308e-18 lub = 1.028216215e-24 wub = 1.403601290e-23 pub = -2.981134876e-30
+ uc = 2.251955405e-10 luc = -3.701600029e-17 wuc = -4.471094413e-16 puc = 8.963416665e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.493074078e-02 lu0 = -9.583780873e-09 wu0 = -1.573237093e-07 pu0 = 3.139159673e-14
+ a0 = 5.123238816e+00 la0 = -9.764893183e-07 wa0 = 1.275264936e-06 pa0 = -2.430654968e-13
+ keta = -1.877737008e-02 lketa = -5.142029332e-09 wketa = 5.707283180e-07 pketa = -1.447545464e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.444921859e+00 lags = 8.977466365e-07 wags = 9.745246929e-07 pags = -2.539611350e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.849812979e-01 lvoff = 1.862417520e-08 wvoff = 7.083140257e-08 pvoff = -1.633985942e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 3.978877490e+00 lnfactor = -1.990423907e-07 wnfactor = -9.915023876e-06 pnfactor = 2.041492786e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.111334796e-05 lcit = -1.593138479e-12 wcit = -1.768988933e-11 pcit = 4.609985160e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -3.020870465e-01 leta0 = 7.790695193e-08 weta0 = 3.308247791e-07 peta0 = -7.766050733e-14
+ etab = -3.582479906e-01 letab = 6.443981004e-08 wetab = 9.528828627e-07 petab = -1.786710207e-13
+ dsub = 8.749634155e-01 ldsub = -1.109972635e-07 wdsub = -2.328895079e-06 pdsub = 4.675090415e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.544024081e+00 lpclm = -2.886626311e-07 wpclm = -2.229423178e-06 ppclm = 5.251687504e-13
+ pdiblc1 = -1.282696956e+00 lpdiblc1 = 4.359048268e-07 wpdiblc1 = 5.742232066e-08 ppdiblc1 = -1.496425676e-14
+ pdiblc2 = 2.474131487e-02 lpdiblc2 = -3.386939267e-09 wpdiblc2 = 1.556526409e-08 ppdiblc2 = -2.015564563e-17
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.734655581e-03 lalpha0 = 8.696587316e-10 walpha0 = 2.237756755e-08 palpha0 = -5.524483637e-15
+ alpha1 = 0.0
+ beta0 = 2.404367742e+01 lbeta0 = 1.692004240e-06 wbeta0 = 3.294175513e-05 pbeta0 = -8.634718900e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 8.962210664e-02 lkt1 = -7.776845691e-08 wkt1 = -7.956698947e-07 pkt1 = 1.604389392e-13
+ kt2 = -1.442438218e-02 lkt2 = -5.792861556e-09 wkt2 = 1.370162094e-08 pkt2 = 1.006270608e-14
+ at = -1.366801920e+05 lat = 4.536918978e-02 wat = 4.479461574e-01 pat = -1.024259522e-7
+ ute = 5.281135183e+00 lute = -1.272068805e-06 wute = -1.992481667e-05 pute = 3.615217379e-12
+ ua1 = 2.108401453e-08 lua1 = -3.876942709e-15 wua1 = -6.067268780e-14 pua1 = 1.114053427e-20
+ ub1 = -1.991916571e-17 lub1 = 3.653306520e-24 wub1 = 5.649458055e-23 pub1 = -1.022593658e-29
+ uc1 = 1.395520365e-10 luc1 = -2.494192275e-17 wuc1 = -6.815233032e-16 puc1 = 1.218076210e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.31 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 2.912482682e-02 lvth0 = 4.216383911e-08 wvth0 = 9.582522211e-07 pvth0 = -1.519873042e-13
+ k1 = 6.328128152e-01 lk1 = 1.660547912e-08 wk1 = 8.566474836e-07 pk1 = -1.784633535e-13
+ k2 = -4.952030899e-02 lk2 = -1.613550659e-08 wk2 = -4.149752653e-07 pk2 = 8.490739304e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.209299539e+05 lvsat = -5.345859952e-03 wvsat = -1.734240469e-01 pvsat = 2.939609521e-8
+ ua = -2.749930259e-09 lua = 1.038028388e-17 wua = 3.298201498e-15 pua = -3.886174584e-22
+ ub = 1.134235365e-18 lub = 3.821505122e-25 wub = 3.723866645e-24 pub = -1.015639799e-30
+ uc = 1.421713030e-10 luc = -2.119158063e-17 wuc = -1.252025730e-16 puc = 2.827871754e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.894861081e-02 lu0 = 6.403623539e-09 wu0 = 1.389197069e-07 pu0 = -2.507239841e-14
+ a0 = 0.0
+ keta = -3.322027448e-01 lketa = 5.459684708e-08 wketa = 1.646032064e-06 pketa = -3.497074405e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.302597604e+00 lags = -7.130573124e-09 wags = -2.106622352e-06 pags = 3.333054917e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = 2.660304154e-01 lvoff = -6.733865735e-08 wvoff = -1.192950639e-06 pvoff = 2.245369976e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.313979636e+00 lnfactor = -2.629128598e-07 wnfactor = -1.063128940e-05 pnfactor = 2.178012994e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.965681037e-05 lcit = -5.127522413e-12 wcit = -1.488015443e-10 pcit = 2.959986660e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.880749005e-01 leta0 = -7.269791517e-08 weta0 = -1.164232341e-06 peta0 = 2.072973797e-13
+ etab = 2.751040814e-02 letab = -9.085740771e-09 wetab = -3.519286268e-07 petab = 7.002604915e-14
+ dsub = 4.671587816e-01 ldsub = -3.326970032e-08 wdsub = 7.873879794e-07 pdsub = -1.264545095e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.031472604e+00 lpclm = 3.928270371e-07 wpclm = 7.160022495e-06 ppclm = -1.264459595e-12
+ pdiblc1 = 2.507556907e+00 lpdiblc1 = -2.865175596e-07 wpdiblc1 = -4.416965545e-06 ppdiblc1 = 8.378540705e-13
+ pdiblc2 = 5.120972761e-02 lpdiblc2 = -8.431818735e-09 wpdiblc2 = -1.216641397e-08 ppdiblc2 = 5.265502192e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.207572646e-02 lalpha0 = -1.762600085e-09 walpha0 = -3.010684210e-08 palpha0 = 4.479044843e-15
+ alpha1 = 0.0
+ beta0 = 4.361902425e+01 lbeta0 = -2.039056867e-06 wbeta0 = -3.269428110e-05 pbeta0 = 3.875509605e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.162162527e+00 lkt1 = 1.608216943e-07 wkt1 = 3.313147246e-06 pkt1 = -6.227016078e-13
+ kt2 = -2.184832330e-01 lkt2 = 3.310075541e-08 wkt2 = 4.112218863e-07 pkt2 = -6.570465650e-14
+ at = 3.433907901e+05 lat = -4.613233941e-02 wat = -1.047623750e+00 pat = 1.826296721e-7
+ ute = -3.088572202e+00 lute = 3.231974223e-07 wute = 3.015374865e-06 pute = -7.571831279e-13
+ ua1 = -9.483701753e-10 lua1 = 3.224298162e-16 wua1 = -8.350988455e-17 pua1 = -4.077630403e-22
+ ub1 = 7.072011298e-19 lub1 = -2.780789993e-25 wub1 = 3.428536872e-24 pub1 = -1.115486532e-31
+ uc1 = 8.917805351e-11 luc1 = -1.534064158e-17 wuc1 = 2.394141033e-16 puc1 = -5.372304865e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.32 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4255045
+ k1 = 0.50407
+ k2 = -0.048314461
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169790.0
+ ua = -1.1014364e-9
+ ub = 2.407218e-18
+ uc = 6.9010287e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0324708
+ a0 = 1.6844032
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5385232
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11480431
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.41179304
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.2558
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.33 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4255045
+ k1 = 0.50407
+ k2 = -0.048314461
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169790.0
+ ua = -1.1014364e-9
+ ub = 2.407218e-18
+ uc = 6.9010287e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0324708
+ a0 = 1.6844032
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5385232
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11480431
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.41179304
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.2558
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.34 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.159485203e-01 lvth0 = 3.832521210e-8
+ k1 = 5.659864270e-01 lk1 = -2.483220221e-7
+ k2 = -7.820229238e-02 lk2 = 1.198681365e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.021648881e+05 lvsat = -5.309027262e-1
+ ua = -9.666125508e-10 lua = -5.407245295e-16
+ ub = 2.261618390e-18 lub = 5.839417943e-25
+ uc = 4.900208962e-11 luc = 8.024487641e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.263164800e-02 lu0 = -6.450969888e-10
+ a0 = 1.546476241e+00 la0 = 5.531698615e-7
+ keta = 2.531445930e-01 lketa = -1.015261705e-6
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.721563730e-01 lags = 4.855551496e-06 pags = 2.067951531e-25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.116893377e-01 lvoff = -1.249290797e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.499306969e+00 lnfactor = -3.509833617e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398762215e-01 letab = 2.802455739e-7
+ dsub = 7.769140535e-01 ldsub = -8.699555029e-07 wdsub = -1.084202172e-19
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.163260720e-01 lpclm = -6.547734436e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 5.433160520e-03 lpdiblc2 = 5.126908318e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.491070895e-05 lalpha0 = 4.160380748e-10 palpha0 = 2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.410270304e+01 lbeta0 = 1.481133413e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.581524020e-01 lkt1 = 9.434543461e-9
+ kt2 = -3.330623020e-02 lkt2 = -5.910701160e-9
+ at = 5.956944909e+05 lat = -1.111796437e+0
+ ute = -1.311968710e+00 lute = 2.044151083e-7
+ ua1 = 1.940438390e-09 lua1 = 5.793777331e-16
+ ub1 = -1.675521700e-18 lub1 = -1.657092890e-24
+ uc1 = -4.012268080e-11 luc1 = -2.686828958e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.35 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.326549068e-01 lvth0 = 4.735351436e-9
+ k1 = 4.472904560e-01 lk1 = -9.671902834e-9
+ k2 = -1.386459694e-02 lk2 = -9.489233912e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.345360400e+03 lvsat = 8.134557942e-2
+ ua = -9.794756888e-10 lua = -5.148619043e-16
+ ub = 2.603000612e-18 lub = -1.024412999e-25
+ uc = 1.044661340e-10 luc = -3.127113122e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.686470711e-02 lu0 = -9.156085626e-9
+ a0 = 2.108717492e+00 la0 = -5.772723972e-7
+ keta = -3.188734160e-01 lketa = 1.348377042e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.429108537e+00 lags = 6.307482667e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.197246989e-01 lvoff = 3.662989369e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 7.287822219e-01 lnfactor = 1.198233694e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.345524140e-04 leta0 = -6.947108359e-11
+ etab = -5.117958520e-04 letab = 3.945973803e-11
+ dsub = -1.014849988e-01 ldsub = 8.961536316e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.784734320e-01 lpclm = -1.904308264e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.682604060e-03 lpdiblc2 = 1.065717714e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.377584428e-04 lalpha0 = -1.925085218e-10
+ alpha1 = 0.0
+ beta0 = 2.213325482e+01 lbeta0 = -1.334893272e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.416056620e-01 lkt1 = -2.383433198e-8
+ kt2 = -5.170615880e-02 lkt2 = 3.108419528e-8
+ at = 7.956296400e+03 lat = 6.990997666e-2
+ ute = -1.315402400e+00 lute = 2.113188854e-7
+ ua1 = 1.752607400e-09 lua1 = 9.570307216e-16
+ ub1 = -1.933764000e-18 lub1 = -1.137870922e-24
+ uc1 = -1.878401720e-11 luc1 = -6.977180662e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.36 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.401908511e-01 lvth0 = -2.880473876e-9
+ k1 = 4.446743720e-01 lk1 = -7.028088343e-9
+ k2 = -1.791730762e-02 lk2 = -5.393564496e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.398586600e+04 lvsat = 1.133214744e-1
+ ua = -1.722316731e-09 lua = 2.358532534e-16
+ ub = 2.906508760e-18 lub = -4.091666343e-25
+ uc = 9.922047680e-11 luc = -2.596987005e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.644243643e-02 lu0 = 1.376661119e-9
+ a0 = 1.262899320e+00 la0 = 2.775114472e-7
+ keta = -3.624720340e-01 lketa = 1.788984676e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.324717717e+00 lags = -1.284954370e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.211672938e-01 lvoff = 5.120875700e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.327511996e+00 lnfactor = 5.931573843e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.312831720e-04 leta0 = -4.704071876e-10
+ etab = -8.540229139e-04 letab = 3.853144068e-10
+ dsub = 5.659857836e-01 ldsub = 2.216076589e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.183971320e-01 lpclm = 2.106465656e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.558901440e-02 lpdiblc2 = -2.386041153e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.642958181e-05 lalpha0 = 6.437389593e-11
+ alpha1 = 0.0
+ beta0 = 1.781694444e+01 lbeta0 = 3.027169998e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.721443720e-01 lkt1 = 7.028088343e-9
+ kt2 = -1.688975120e-02 lkt2 = -4.101266237e-9
+ at = 8.251676640e+04 lat = -5.440834324e-3
+ ute = -6.610568000e-01 lute = -4.499627779e-7
+ ua1 = 5.155208156e-09 lua1 = -2.481637602e-15
+ ub1 = -6.116866440e-18 lub1 = 3.089572404e-24
+ uc1 = -1.775098688e-10 luc1 = 9.063653901e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.37 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.006786576e-01 lvth0 = -3.376554787e-8
+ k1 = 2.648519899e-01 lk1 = 8.478921996e-8
+ k2 = 2.687543262e-02 lk2 = -2.826473766e-08 pk2 = -1.615587134e-27
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.928791329e+05 lvsat = -2.515794073e-3
+ ua = -1.994271278e-10 lua = -5.417341782e-16
+ ub = 1.602399052e-18 lub = 2.567117822e-25
+ uc = 4.924934511e-11 luc = -4.546102142e-19
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.344405666e-02 lu0 = -7.304366173e-9
+ a0 = 2.131485262e+00 la0 = -1.659885345e-7
+ keta = 9.924730893e-03 lketa = -1.124732059e-08 pketa = 8.077935669e-28
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.650585984e+00 lags = -4.301427074e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.115896756e-01 lvoff = 2.305438449e-10
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.482255469e+00 lnfactor = 3.545366745e-9
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -8.534188585e-03 leta0 = 4.362662692e-09 weta0 = -2.911675756e-22 peta0 = 1.443615457e-28
+ etab = 1.919533138e-02 letab = -9.851885895e-09 wetab = -3.705769144e-22 petab = 4.985600921e-28
+ dsub = 1.767026398e+00 ldsub = -3.916436790e-07 wdsub = -2.168404345e-19 pdsub = 5.169878828e-26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.230923648e-01 lpclm = 3.628202854e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.472925600e-03 lpdiblc2 = 3.289833789e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.871020363e-03 lalpha0 = 1.011327949e-09 walpha0 = -2.646977960e-23 palpha0 = 2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.673611267e+01 lbeta0 = 3.579042699e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.452144880e-01 lkt1 = -6.722310427e-9
+ kt2 = -3.153915520e-02 lkt2 = 3.378719445e-9
+ at = 8.798797040e+04 lat = -8.234431086e-3
+ ute = -1.386565440e+00 lute = -7.951806634e-8
+ ua1 = 5.888173480e-10 lua1 = -1.500384559e-16
+ ub1 = -2.000359616e-19 lub1 = 6.843876199e-26 pub1 = 5.605193857e-45
+ uc1 = 3.142940240e-11 luc1 = -1.604785287e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.38 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.486027986e-01 lvth0 = -4.625457901e-8
+ k1 = 3.119744075e-01 lk1 = 7.250911793e-8
+ k2 = 3.291655585e-02 lk2 = -2.983905438e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.749921224e+05 lvsat = 2.145560871e-3
+ ua = -2.327078853e-09 lua = 1.273186146e-17
+ ub = 2.595219338e-18 lub = -2.017184277e-27
+ uc = 7.068153865e-11 luc = -6.039839851e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.056213734e-02 lu0 = 1.264662003e-9
+ a0 = 5.563950352e+00 la0 = -1.060488937e-6
+ keta = 1.784573743e-01 lketa = -5.516692745e-08 wketa = 1.355252716e-20 pketa = -3.231174268e-27
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.108141429e+00 lags = 8.099816563e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.605030774e-01 lvoff = 1.297737638e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 5.524009374e-01 lnfactor = 5.064654578e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.877591979e-01 leta0 = 5.106870013e-08 weta0 = -3.388131789e-21 peta0 = -2.423380701e-27
+ etab = -2.894663676e-02 letab = 2.693911001e-9
+ dsub = 7.013384757e-02 ldsub = 5.056651973e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 7.735704401e-01 lpclm = -1.071725579e-7
+ pdiblc1 = -1.262852704e+00 lpdiblc1 = 4.307334147e-7
+ pdiblc2 = 3.012042571e-02 lpdiblc2 = -3.393904741e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.998680363e-03 lalpha0 = -1.039516060e-9
+ alpha1 = 0.0
+ beta0 = 3.542783069e+01 lbeta0 = -1.292019018e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.853489143e-01 lkt1 = -2.232327894e-8
+ kt2 = -9.689317143e-03 lkt2 = -2.315348353e-9
+ at = 1.812296571e+04 lat = 9.972389135e-3
+ ute = -1.604568571e+00 lute = -2.270645029e-8
+ ua1 = 1.164863914e-10 lua1 = -2.694900861e-17 wua1 = 6.310887242e-30 pua1 = -1.504632769e-36
+ ub1 = -3.955258229e-19 lub1 = 1.193834198e-25
+ uc1 = -9.597171486e-11 luc1 = 1.715287829e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.39 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.018908126e+00 lvth0 = 6.337130033e-07 wvth0 = 9.778192776e-06 pvth0 = -1.863723543e-12
+ k1 = 9.288567333e-01 lk1 = -4.506865337e-8
+ k2 = 9.463316632e-01 lk2 = -2.039359738e-07 wk2 = -3.296622325e-06 pk2 = 6.283362151e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.272560921e+06 lvsat = -1.160051052e+00 wvsat = -1.768472599e+01 pvsat = 3.370708774e-6
+ ua = -8.710916099e-09 lua = 1.229491240e-15 wua = 2.054720817e-14 pua = -3.916297878e-21
+ ub = 2.688314546e-17 lub = -4.631295903e-24 wub = -7.078446705e-23 pub = 1.349151942e-29
+ uc = 9.890325989e-11 luc = -1.141889992e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -9.967044928e-02 lu0 = 2.227499301e-08 wu0 = 3.725004548e-07 pu0 = -7.099858669e-14
+ a0 = 0.0
+ keta = 2.366400884e-01 lketa = -6.625655277e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.745820000e-01 lags = 1.080545708e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.462345920e-01 lvoff = 1.025780305e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -7.839818213e+01 lnfactor = 1.555444659e-05 wnfactor = 2.287087575e-04 pnfactor = -4.359188918e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 8.573448585e-02 leta0 = -1.059196002e-9
+ etab = -9.411059882e-02 letab = 1.511416217e-8
+ dsub = 7.392677026e-01 ldsub = -7.697039304e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.429187333e-01 lpclm = -4.415034257e-8
+ pdiblc1 = 9.811229760e-01 lpdiblc1 = 3.031650054e-9
+ pdiblc2 = 4.700520600e-02 lpdiblc2 = -6.612143864e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.671274608e-03 lalpha0 = -2.147125235e-10
+ alpha1 = 0.0
+ beta0 = 3.232039411e+01 lbeta0 = -6.997416058e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.719086667e-02 lkt1 = -5.437420281e-8
+ kt2 = -7.637140667e-02 lkt2 = 1.039425791e-8
+ at = -1.865152667e+04 lat = 1.698160738e-2
+ ute = -2.046506000e+00 lute = 6.152682360e-8
+ ua1 = -9.772298800e-10 lua1 = 1.815133127e-16 wua1 = 2.524354897e-29 pua1 = -6.018531076e-36
+ ub1 = 1.892049633e-18 lub1 = -3.166284621e-25 wub1 = 1.880790961e-37 pub1 = 2.242077543e-44
+ uc1 = 1.719158080e-10 luc1 = -3.390648356e-17 wuc1 = 6.310887242e-30 puc1 = 2.256949154e-36
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.40 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.300018434e-01 wvth0 = -1.296876436e-8
+ k1 = 4.709090789e-01 wk1 = 9.562449016e-8
+ k2 = -3.781288124e-02 wk2 = -3.028288049e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.348455007e+05 wvsat = 1.007677053e-1
+ ua = -1.240718153e-09 wua = 4.016398280e-16
+ ub = 2.717296924e-18 wub = -8.941590880e-25
+ uc = 1.220174343e-10 wuc = -1.528540604e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.620449933e-02 wu0 = -1.076668206e-8
+ a0 = 1.421338942e+00 wa0 = 7.585852476e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.957823058e-01 wags = 1.232497797e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.199962492e-01 wvoff = 1.497173544e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 9.409661708e-01 wnfactor = 1.357699901e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.801851852e-07 wcit = 1.637966601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 5.737234637e-03 wpdiblc2 = 2.809440314e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.551688192e-05 walpha0 = 9.536320173e-12
+ alpha1 = 0.0
+ beta0 = 1.779846172e+01 wbeta0 = -7.819652553e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.537210522e-01 wkt1 = -5.994957759e-9
+ kt2 = -3.298051733e-02 wkt2 = -5.189078192e-9
+ at = 6.141336389e+05 wat = -8.525616158e-1
+ ute = -1.352110170e+00 wute = 2.627298428e-7
+ ua1 = 2.222701293e-09 wua1 = -3.973706974e-16
+ ub1 = -2.796110263e-18 wub1 = 2.039923605e-24
+ uc1 = -1.720587230e-10 wuc1 = 3.611388762e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.41 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.300018434e-01 wvth0 = -1.296876436e-8
+ k1 = 4.709090789e-01 wk1 = 9.562449016e-8
+ k2 = -3.781288124e-02 wk2 = -3.028288049e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.348455007e+05 wvsat = 1.007677053e-1
+ ua = -1.240718153e-09 wua = 4.016398280e-16
+ ub = 2.717296924e-18 wub = -8.941590880e-25
+ uc = 1.220174343e-10 wuc = -1.528540604e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.620449933e-02 wu0 = -1.076668206e-8
+ a0 = 1.421338942e+00 wa0 = 7.585852476e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.957823058e-01 wags = 1.232497797e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.199962492e-01 wvoff = 1.497173544e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 9.409661708e-01 wnfactor = 1.357699901e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.801851852e-07 wcit = 1.637966601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 5.737234637e-03 wpdiblc2 = 2.809440314e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.551688192e-05 walpha0 = 9.536320173e-12
+ alpha1 = 0.0
+ beta0 = 1.779846172e+01 wbeta0 = -7.819652553e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.537210522e-01 wkt1 = -5.994957759e-9
+ kt2 = -3.298051733e-02 wkt2 = -5.189078192e-9
+ at = 6.141336389e+05 wat = -8.525616158e-1
+ ute = -1.352110170e+00 wute = 2.627298428e-7
+ ua1 = 2.222701293e-09 wua1 = -3.973706974e-16
+ ub1 = -2.796110263e-18 wub1 = 2.039923605e-24
+ uc1 = -1.720587230e-10 wuc1 = 3.611388762e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.42 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.274691780e-01 lvth0 = 1.015750782e-08 wvth0 = -3.322154460e-08 pvth0 = 8.122580045e-14
+ k1 = 5.171336285e-01 lk1 = -1.853881787e-07 wk1 = 1.408743724e-07 pk1 = -1.814791776e-13
+ k2 = -6.818409211e-02 lk2 = 1.218067783e-07 wk2 = -2.888898322e-08 pk2 = -5.590364362e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.373270198e+05 lvsat = -4.110123804e-01 wvsat = 1.869697189e-01 pvsat = -3.457217957e-7
+ ua = -1.099315171e-09 lua = -5.671108029e-16 wua = 3.826679092e-16 pua = 7.608877742e-23
+ ub = 2.576465292e-18 lub = 5.648193414e-25 wub = -9.079082680e-25 pub = 5.514246131e-32
+ uc = 1.125295329e-10 luc = 3.805217733e-17 wuc = -1.831909119e-16 puc = 1.216689767e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.670739371e-02 lu0 = -2.016908204e-09 wu0 = -1.175302411e-08 pu0 = 3.955823412e-15
+ a0 = 1.047262819e+00 la0 = 1.500269699e-06 wa0 = 1.439556785e-06 pa0 = -2.731104446e-12
+ keta = 3.337510490e-01 lketa = -1.338541957e-06 wketa = -2.324408068e-07 pketa = 9.322270998e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -1.104604928e+00 lags = 6.418513039e-06 wags = 1.247030275e-06 pags = -4.507034054e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.211150345e-01 lvoff = 4.487000252e-09 wvoff = 2.718041053e-08 pvoff = -4.896411234e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 5.147423325e-01 lnfactor = 1.709413326e-06 wnfactor = 2.839139813e-06 pnfactor = -5.941462908e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.801851852e-07 wcit = 1.637966601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398851638e-01 letab = 2.802814380e-07 wetab = 2.578650492e-11 petab = -1.034193566e-16
+ dsub = 8.431688943e-01 ldsub = -1.135677168e-06 wdsub = -1.910557717e-07 pdsub = 7.662482781e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.743083584e-01 lpclm = -2.980211020e-07 wpclm = -1.672006200e-07 ppclm = 6.705748067e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 7.779200477e-03 lpdiblc2 = -8.189508199e-09 wpdiblc2 = -6.765158123e-09 ppdiblc2 = 3.839988449e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.161597834e-05 lalpha0 = 5.098790493e-10 walpha0 = 7.700865005e-11 palpha0 = -2.706045262e-16
+ alpha1 = 0.0
+ beta0 = 1.379054365e+01 lbeta0 = 1.607415620e-05 wbeta0 = 9.001584240e-07 pbeta0 = -3.641536874e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.711828820e-01 lkt1 = 7.003241452e-08 wkt1 = 3.757534366e-08 pkt1 = -1.747430509e-13
+ kt2 = -3.066048253e-02 lkt2 = -9.304731580e-09 wkt2 = -7.629410267e-09 pkt2 = 9.787195820e-15
+ at = 1.195929297e+06 lat = -2.333349666e+00 wat = -1.730867099e+00 pat = 3.522531969e-6
+ ute = -1.391201477e+00 lute = 1.567795937e-07 wute = 2.284795681e-07 pute = 1.373641519e-13
+ ua1 = 2.008574143e-09 lua1 = 8.587783479e-16 wua1 = -1.964796629e-16 pua1 = -8.056935830e-22
+ ub1 = -2.402689567e-18 lub1 = -1.577853043e-24 wub1 = 2.096897620e-24 pub1 = -2.284999834e-31
+ uc1 = -2.406713929e-10 luc1 = 2.751779741e-16 wuc1 = 5.783122937e-16 puc1 = -8.709957083e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.43 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.331664104e-01 lvth0 = -1.297347584e-09 wvth0 = -1.474997343e-09 pvth0 = 1.739619253e-14
+ k1 = 4.346869044e-01 lk1 = -1.962079521e-08 wk1 = 3.634423158e-08 pk1 = 2.868912349e-14
+ k2 = -2.014123538e-03 lk2 = -1.123456048e-08 wk2 = -3.417261763e-08 pk2 = 5.032910968e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -5.988110418e+03 lvsat = 7.819702044e-02 wvsat = 1.050441609e-02 pvsat = 9.079342099e-9
+ ua = -1.298002379e-09 lua = -1.676303024e-16 wua = 9.185194890e-16 pua = -1.001294409e-21
+ ub = 3.021893421e-18 lub = -3.307584541e-25 wub = -1.207940249e-24 pub = 6.583867616e-31
+ uc = 1.567189014e-10 luc = -5.079496688e-17 wuc = -1.506786927e-16 puc = 5.629990870e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.968348320e-02 lu0 = -8.000633730e-09 wu0 = -8.128363673e-09 pu0 = -3.331918858e-15
+ a0 = 2.001871513e+00 la0 = -4.190665418e-07 wa0 = 3.081064060e-07 pa0 = -4.562103148e-13
+ keta = -3.963454436e-01 lketa = 1.293900508e-07 wketa = 2.234022123e-07 pketa = 1.570912563e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.761241475e+00 lags = 6.564422623e-07 wags = -9.577551442e-07 pags = -7.409249040e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.206054905e-01 lvoff = 3.462511108e-09 wvoff = 2.539894532e-09 pvoff = 5.781091358e-16
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.003696977e+00 lnfactor = 7.263211185e-07 wnfactor = -7.927579322e-07 pnfactor = 1.360830698e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.420580333e-06 lcit = 1.154163848e-11 wcit = 3.293295648e-11 pcit = -3.328204582e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.974350190e-04 leta0 = 5.157150855e-12 weta0 = 1.070335762e-10 peta0 = -2.152017083e-16
+ etab = -4.929468368e-04 letab = 1.944653690e-11 wetab = -5.435396264e-11 petab = 5.771106745e-17
+ dsub = -4.780043780e-01 ldsub = 1.520673814e-06 wdsub = 1.085750108e-06 pdsub = -1.800897623e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.024367314e-01 lpclm = -3.545760089e-07 wpclm = -6.910176839e-08 ppclm = 4.733372556e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -4.234928741e-03 lpdiblc2 = 1.596610001e-08 wpdiblc2 = 1.994774346e-08 ppdiblc2 = -1.530907543e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.776641528e-04 lalpha0 = -2.325955823e-10 walpha0 = -1.150741005e-10 palpha0 = 1.155970520e-16
+ alpha1 = 0.0
+ beta0 = 2.272318965e+01 lbeta0 = -1.885821843e-06 wbeta0 = -1.701165583e-06 pbeta0 = 1.588685175e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.121895370e-01 lkt1 = -4.857960489e-08 wkt1 = -8.482580879e-08 pkt1 = 7.135670623e-14
+ kt2 = -5.180815652e-02 lkt2 = 3.321478175e-08 wkt2 = 2.941257314e-10 pkt2 = -6.143865658e-15
+ at = -5.134559428e+03 lat = 8.150932334e-02 wat = 3.774944641e-02 pat = -3.344845605e-8
+ ute = -1.506959057e+00 lute = 3.895217836e-07 wute = 5.523823529e-07 pute = -5.138747874e-13
+ ua1 = 1.360754122e-09 lua1 = 2.161285281e-15 wua1 = 1.129967705e-15 pua1 = -3.472648661e-21
+ ub1 = -1.784915633e-18 lub1 = -2.819949314e-24 wub1 = -4.292265925e-25 pub1 = 4.850525357e-30
+ uc1 = -7.648668546e-11 luc1 = -5.493179869e-17 wuc1 = 1.663942993e-16 puc1 = -4.279338887e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.44 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.296327147e-01 lvth0 = 2.273805270e-09 wvth0 = 3.044596999e-08 pvth0 = -1.486313706e-14
+ k1 = 4.480041693e-01 lk1 = -3.307922308e-08 wk1 = -9.601969874e-09 pk1 = 7.512235469e-14
+ k2 = -1.005872965e-02 lk2 = -3.104681549e-09 wk2 = -2.266138838e-08 pk2 = -6.600337309e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.604682031e+04 lvsat = 1.085743527e-01 wvsat = 5.943070909e-03 pvsat = 1.368903754e-8
+ ua = -2.361542113e-09 lua = 9.071829528e-16 wua = 1.843302270e-15 pua = -1.935879888e-21
+ ub = 3.627576490e-18 lub = -9.428617641e-25 wub = -2.079306961e-24 pub = 1.538989961e-30
+ uc = 1.755322420e-10 luc = -6.980772890e-17 wuc = -2.200564217e-16 puc = 1.264130417e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.514450765e-02 lu0 = 6.692454956e-09 wu0 = 3.742772324e-09 pu0 = -1.532888890e-14
+ a0 = 4.024488986e-01 la0 = 1.197309952e-06 wa0 = 2.481237858e-06 pa0 = -2.652376960e-12
+ keta = -5.159129463e-01 lketa = 2.502249691e-07 wketa = 4.424698867e-07 pketa = -2.056806661e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.372605206e+00 lags = -9.720019247e-07 wags = -1.380907569e-07 pags = -9.024453202e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.369106805e-01 lvoff = 1.994053618e-08 wvoff = 4.539841727e-08 pvoff = -4.273471394e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 3.509115586e-01 lnfactor = 1.386026062e-06 wnfactor = 2.816173851e-06 pnfactor = -2.286355762e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.138029529e-03 leta0 = -3.674027661e-09 weta0 = -9.247134133e-09 peta0 = 9.238120179e-15
+ etab = -8.856597526e-04 letab = 4.163222095e-10 wetab = 9.122956984e-11 petab = -8.941565048e-17
+ dsub = 1.054005179e+00 ldsub = -2.757504423e-08 wdsub = -1.407277128e-06 pdsub = 7.185557018e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.626371609e-01 lpclm = 3.175476667e-07 wpclm = 7.043027593e-07 ppclm = -3.082653601e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 8.083046745e-03 lpdiblc2 = 3.517553981e-09 wpdiblc2 = 2.164458363e-08 ppdiblc2 = -1.702390211e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.024104834e-05 lalpha0 = 2.755620706e-11 walpha0 = -1.057452626e-10 palpha0 = 1.061693285e-16
+ alpha1 = 0.0
+ beta0 = 1.853258551e+01 lbeta0 = 2.349202699e-06 wbeta0 = -2.063658386e-06 pbeta0 = 1.955020401e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.764485346e-01 lkt1 = 1.636053805e-08 wkt1 = 1.241169847e-08 pkt1 = -2.691151860e-14
+ kt2 = -2.545105218e-02 lkt2 = 6.578292103e-09 wkt2 = 2.468779558e-08 pkt2 = -3.079610841e-14
+ at = 9.031797590e+04 lat = -1.495500887e-02 wat = -2.249595778e-02 pat = 2.743554943e-8
+ ute = -2.125793237e-01 lute = -9.185783745e-07 wute = -1.293252074e-06 pute = 1.351323365e-12
+ ua1 = 8.124323333e-09 lua1 = -4.673977764e-15 wua1 = -8.561888981e-15 pua1 = 6.321941706e-21
+ ub1 = -1.060259529e-17 lub1 = 6.091197749e-24 wub1 = 1.293527200e-23 pub1 = -8.655636925e-30
+ uc1 = -2.780388627e-10 luc1 = 1.487568316e-16 wuc1 = 2.898904333e-16 puc1 = -1.675985819e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.45 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.909045710e-01 lvth0 = -2.901160454e-08 wvth0 = 2.818504486e-08 pvth0 = -1.370870869e-14
+ k1 = 1.796413484e-01 lk1 = 1.039468333e-07 wk1 = 2.457176665e-07 pk1 = -5.524385163e-14
+ k2 = 5.994307163e-02 lk2 = -3.884760128e-08 wk2 = -9.535549725e-08 pk2 = 3.051727468e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.406173147e+05 lvsat = 1.836964531e-02 wvsat = 1.507047920e-01 pvsat = -6.022629727e-8
+ ua = 1.255936096e-09 lua = -9.399014207e-16 wua = -4.196758162e-15 pua = 1.148174969e-21
+ ub = 4.733019163e-19 lub = 6.677108333e-25 wub = 3.255920957e-24 pub = -1.185177414e-30
+ uc = 2.303437926e-11 luc = 8.057679817e-18 wuc = 7.559478627e-17 puc = -2.454646515e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.858375227e-02 lu0 = -1.038162335e-08 wu0 = -4.365758324e-08 pu0 = 8.873732653e-15
+ a0 = 4.077171639e+00 la0 = -6.790034786e-07 wa0 = -5.610678522e-06 pa0 = 1.479355543e-12
+ keta = -1.089994895e-02 lketa = -7.634667343e-09 wketa = 6.005108802e-08 pketa = -1.041762753e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.000201174e+00 lags = -7.818524259e-07 wags = -3.891817843e-06 pags = 1.014207730e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -8.555414408e-02 lvoff = -6.282111335e-09 wvoff = -7.507736035e-08 pvoff = 1.878021811e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 3.237936554e+00 lnfactor = -8.808890083e-08 wnfactor = -2.179119760e-06 pnfactor = 2.642411557e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.092102504e-05 lcit = -3.023275384e-12 wcit = -1.707416385e-11 pcit = 8.718068061e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.112008228e-02 leta0 = 9.222764226e-09 weta0 = 3.629331234e-08 peta0 = -1.401483179e-14
+ etab = 3.109951072e-02 letab = -1.591530583e-08 wetab = -3.432748675e-08 petab = 1.748478090e-14
+ dsub = 1.867905010e+00 ldsub = -4.431522980e-07 wdsub = -2.908986079e-07 pdsub = 1.485328292e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.845129998e-01 lpclm = -6.394720537e-08 wpclm = -4.654806140e-07 ppclm = 2.890260304e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 7.094249450e-03 lpdiblc2 = 4.022433880e-09 wpdiblc2 = -7.558980520e-09 ppdiblc2 = -2.112562252e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.646910139e-03 lalpha0 = 1.389403603e-09 walpha0 = 2.237394554e-09 palpha0 = -1.090237862e-15
+ alpha1 = 0.0
+ beta0 = 1.484878072e+01 lbeta0 = 4.230153425e-06 wbeta0 = 5.442404770e-06 pbeta0 = -1.877575446e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.169360360e-01 lkt1 = -1.402654375e-08 wkt1 = -8.154515824e-08 pkt1 = 2.106285243e-14
+ kt2 = -1.330754297e-02 lkt2 = 3.778162990e-10 wkt2 = -5.257358861e-08 pkt2 = 8.653554357e-15
+ at = 6.201579623e+04 lat = -5.039159296e-04 wat = 7.489466004e-02 pat = -2.229210003e-8
+ ute = -1.549745346e+00 lute = -2.358214037e-07 wute = 4.705537347e-07 pute = 4.507241187e-13
+ ua1 = -7.840437999e-10 lua1 = -1.253655055e-16 wua1 = 3.958851049e-15 pua1 = -7.114815344e-23
+ ub1 = 1.553314475e-18 lub1 = -1.156097782e-25 wub1 = -5.056048986e-24 pub1 = 5.307315730e-31
+ uc1 = 1.028517127e-10 luc1 = -4.572589614e-17 wuc1 = -2.059569450e-16 puc1 = 8.558108948e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.46 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.564652574e-01 lvth0 = -4.609671942e-08 wvth0 = -2.267257935e-08 pvth0 = -4.552118188e-16
+ k1 = 3.856932875e-01 lk1 = 5.024969793e-08 wk1 = -2.125794483e-07 pk1 = 6.418837648e-14
+ k2 = -8.770342405e-03 lk2 = -2.094088558e-08 wk2 = 1.202104242e-07 pk2 = -2.565920444e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.852664659e+05 lvsat = -1.932592348e-02 wvsat = -3.179926105e-01 pvsat = 6.191624584e-8
+ ua = -2.630988136e-09 lua = 7.303103427e-17 wua = 8.763680030e-16 pua = -1.738817097e-22
+ ub = 3.492522958e-18 lub = -1.190981702e-25 wub = -2.587509583e-24 pub = 3.376205850e-31
+ uc = 6.952147748e-11 luc = -4.056857978e-18 wuc = 3.345210410e-18 puc = -5.718225678e-24
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.664838189e-02 lu0 = 5.467341739e-10 wu0 = -1.755059909e-08 pu0 = 2.070252584e-15
+ a0 = 5.478677864e+00 la0 = -1.044236001e-06 wa0 = 2.458960098e-07 pa0 = -4.686777947e-14
+ keta = 1.775565937e-01 lketa = -5.674644235e-08 wketa = 2.597535920e-09 pketa = 4.554768147e-15
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.253524957e+00 lags = 8.478686038e-07 wags = 4.192352116e-07 pags = -1.092526961e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.429053962e-01 lvoff = 8.663624962e-09 wvoff = -5.074555358e-08 pvoff = 1.243934926e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.358253406e+00 lnfactor = 1.411565275e-07 wnfactor = -5.207446472e-06 pnfactor = 1.053423097e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.614651799e-05 lcit = 4.030526329e-12 wcit = 6.097915660e-11 pcit = -1.162262725e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.831542407e-01 leta0 = 5.144886590e-08 weta0 = -1.327908505e-08 peta0 = -1.096265031e-15
+ etab = -8.724984675e-02 letab = 1.492653672e-08 wetab = 1.681260515e-07 petab = -3.527461117e-14
+ dsub = -2.794295123e-01 ldsub = 1.164430784e-07 wdsub = 1.008018383e-06 pdsub = -1.899649385e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.224245586e-02 lpclm = 2.524849837e-08 wpclm = 2.108893942e-06 ppclm = -3.818559788e-13
+ pdiblc1 = -1.253661990e+00 lpdiblc1 = 4.283383147e-07 wpdiblc1 = -2.650280129e-08 ppdiblc1 = 6.906630016e-15
+ pdiblc2 = 5.680678936e-02 lpdiblc2 = -8.932654022e-09 wpdiblc2 = -7.695413254e-08 ppdiblc2 = 1.597181436e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.286584906e-03 lalpha0 = -1.459865205e-09 walpha0 = -6.597515935e-09 palpha0 = 1.212139812e-15
+ alpha1 = 0.0
+ beta0 = 3.675506836e+01 lbeta0 = -1.478625132e-06 wbeta0 = -3.827288887e-06 pbeta0 = 5.381067209e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.897079533e-01 lkt1 = -2.112218209e-08 wkt1 = 1.256994289e-08 pkt1 = -3.463542920e-15
+ kt2 = 1.834263369e-02 lkt2 = -7.870219739e-09 wkt2 = -8.083433502e-08 pkt2 = 1.601830487e-14
+ at = 4.297921589e+04 lat = 4.457016907e-03 wat = -7.167672583e-02 pat = 1.590440313e-8
+ ute = -4.555707811e+00 lute = 5.475324147e-07 wute = 8.510052667e-06 pute = -1.644369303e-12
+ ua1 = -5.302841914e-09 lua1 = 1.052233283e-15 wua1 = 1.562744607e-14 pua1 = -3.111984015e-21
+ ub1 = 4.158888082e-18 lub1 = -7.946222602e-25 wub1 = -1.313333566e-23 pub1 = 2.635672479e-30
+ uc1 = -2.025037471e-10 luc1 = 3.384973666e-17 wuc1 = 3.072010946e-16 puc1 = -4.814789564e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.47 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 6.364032786e-01 lvth0 = -6.133290625e-08 wvth0 = -7.624459567e-07 pvth0 = 1.405455939e-13
+ k1 = 6.552366842e-01 lk1 = -1.125273490e-09 wk1 = 7.890244545e-07 pk1 = -1.267173274e-13
+ k2 = -1.283558755e-01 lk2 = 1.852117018e-09 wk2 = -1.975996037e-07 pk2 = 3.491538688e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.284493351e+05 lvsat = 1.056342164e-02 wvsat = 3.274137990e-02 pvsat = -4.933652737e-9
+ ua = -1.472883926e-09 lua = -1.477036282e-16 wua = -3.247433018e-16 pua = 5.505010503e-23
+ ub = 3.354447214e-18 lub = -9.278093336e-26 wub = -2.935936356e-24 pub = 4.040307277e-31
+ uc = 1.576324003e-10 luc = -2.085079987e-17 wuc = -1.693542858e-16 puc = 2.719829830e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.020213322e-02 lu0 = -3.942610829e-09 wu0 = -3.084311770e-08 pu0 = 4.603806631e-15
+ a0 = 0.0
+ keta = 1.782666324e-01 lketa = -5.688177573e-08 wketa = 1.683286164e-07 pketa = -2.703357580e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.138102328e-01 lags = 5.357451661e-08 wags = -9.782154936e-07 pags = 1.571014083e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.782223708e-01 lvoff = 1.539504033e-08 wvoff = 9.224155843e-08 pvoff = -1.481399428e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -2.025308647e+00 lnfactor = 9.766634548e-07 wnfactor = 8.476120878e-06 pnfactor = -1.554664840e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.276635068e-01 leta0 = -7.792996772e-09 weta0 = -1.209086214e-07 peta0 = 1.941792459e-14
+ etab = -5.677613555e-02 letab = 9.118247369e-09 wetab = -1.076595250e-07 petab = 1.729011972e-14
+ dsub = 7.142604469e-01 ldsub = -7.295422777e-08 wdsub = 7.211217301e-08 pdsub = -1.158121499e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.105834819e-01 lpclm = -6.837301201e-09 wpclm = 6.699735477e-07 ppclm = -1.075977518e-13
+ pdiblc1 = 9.596779776e-01 lpdiblc1 = 6.475716800e-09 wpdiblc1 = 6.183986967e-08 ppdiblc1 = -9.931483070e-15
+ pdiblc2 = 3.192759369e-02 lpdiblc2 = -4.190679327e-09 wpdiblc2 = 4.347855673e-08 ppdiblc2 = -6.982656210e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.195456641e-03 lalpha0 = -2.988961581e-10 walpha0 = -1.511557521e-09 palpha0 = 2.427561378e-16
+ alpha1 = 0.0
+ beta0 = 3.453257360e+01 lbeta0 = -1.055017631e-06 wbeta0 = -6.379151365e-06 pbeta0 = 1.024491709e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.848733089e-03 lkt1 = -5.635634947e-08 wkt1 = -3.559039349e-08 pkt1 = 5.715817195e-15
+ kt2 = -8.343745858e-02 lkt2 = 1.152906585e-08 wkt2 = 2.037602060e-08 pkt2 = -3.272388909e-15
+ at = -4.457722480e+04 lat = 2.114527450e-02 wat = 7.476063943e-02 pat = -1.200655869e-8
+ ute = -1.788115133e+00 lute = 2.002925041e-08 wute = -7.451088228e-07 pute = 1.196644769e-13
+ ua1 = 5.647140083e-10 lua1 = -6.612287574e-17 wua1 = -4.446426494e-15 pua1 = 7.140960949e-22
+ ub1 = 3.609033075e-19 lub1 = -7.072636218e-26 wub1 = 4.415290103e-24 pub1 = -7.090955905e-31
+ uc1 = 5.164424245e-11 luc1 = -1.459087014e-17 wuc1 = 3.468211000e-16 puc1 = -5.569946866e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.48 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.49 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.50 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.058074269e-01 lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-1
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16 puc = 2.350988702e-38
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.033923399e-01 lvoff = -2.743952297e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.365972934e+00 lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10 palpha0 = 4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095730e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.51 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.322046542e-01 lvth0 = 1.004565279e-8
+ k1 = 4.583847700e-01 lk1 = -9.143605620e-10
+ k2 = -2.429601160e-02 lk2 = -7.952904977e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.611812000e+02 lvsat = 8.411710788e-2
+ ua = -6.990916173e-10 lua = -8.205135605e-16
+ ub = 2.234268964e-18 lub = 9.853555799e-26
+ uc = 5.847047920e-11 luc = -1.408521648e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.438347102e-02 lu0 = -1.017317561e-8
+ a0 = 2.202768984e+00 la0 = -7.165335746e-7
+ keta = -2.506784320e-01 lketa = 1.396330174e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.136747526e+00 lags = 6.081310502e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.189493795e-01 lvoff = 3.839460957e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.867876868e-01 lnfactor = 1.613636150e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.672251120e-04 leta0 = -1.351628102e-10
+ etab = -5.283877540e-04 letab = 5.707641819e-11
+ dsub = 2.299473109e-01 ldsub = 3.464178733e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.573796660e-01 lpclm = -4.594153846e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.771783000e-03 lpdiblc2 = 5.983981900e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.026313223e-04 lalpha0 = -1.572217669e-10
+ alpha1 = 0.0
+ beta0 = 2.161396292e+01 lbeta0 = -8.499367487e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.674992940e-01 lkt1 = -2.052231484e-9
+ kt2 = -5.161637500e-02 lkt2 = 2.920874017e-8
+ at = 1.947956140e+04 lat = 5.969961705e-2
+ ute = -1.146784080e+00 lute = 5.445525125e-8
+ ua1 = 2.097537420e-09 lua1 = -1.030179567e-16
+ ub1 = -2.064788220e-18 lub1 = 3.427836151e-25
+ uc1 = 3.200892914e-11 luc1 = -8.283476799e-17 wuc1 = -6.162975822e-33
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.52 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.494846822e-01 lvth0 = -7.417543512e-9
+ k1 = 4.417433080e-01 lk1 = 1.590350094e-8
+ k2 = -2.483484439e-02 lk2 = -7.408360556e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.217170480e+04 lvsat = 1.175001425e-01 pvsat = 2.646977960e-23
+ ua = -1.159636678e-09 lua = -3.550867226e-16
+ ub = 2.271786733e-18 lub = 6.062010003e-26
+ uc = 3.204681721e-11 luc = 1.261853632e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.758494212e-02 lu0 = -3.302582306e-9
+ a0 = 2.020313377e+00 la0 = -5.321439384e-7
+ keta = -2.274052120e-01 lketa = 1.161131012e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.282564612e+00 lags = -1.560431697e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.073091305e-01 lvoff = -7.924174767e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.187167452e+00 lnfactor = -1.047676407e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.891464901e-03 leta0 = 2.349589317e-09 weta0 = 4.135903063e-25 peta0 = -1.972152263e-31
+ etab = -8.261744920e-04 letab = 3.580196956e-10
+ dsub = 1.364052514e-01 ldsub = 4.409514786e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.659588400e-02 lpclm = 1.165465516e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.219616488e-02 lpdiblc2 = -7.582698428e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.870901370e-05 lalpha0 = 9.678277668e-11 palpha0 = -1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.718699924e+01 lbeta0 = 3.623952740e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.683556200e-01 lkt1 = -1.186828428e-9
+ kt2 = -9.353640400e-03 lkt2 = -1.350197941e-8
+ at = 7.564972840e+04 lat = 2.934046279e-3
+ ute = -1.055830440e+00 lute = -3.746249734e-8
+ ua1 = 2.541635640e-09 lua1 = -5.518236178e-16
+ ub1 = -2.168290200e-18 lub1 = 4.473827161e-25
+ uc1 = -8.901892120e-11 luc1 = 3.947597756e-17 wuc1 = 2.465190329e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.53 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.092823266e-01 lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.345075300e-01 lvoff = 5.963328048e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.817064934e+00 lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 7.237830360e-25 petab = -3.451266460e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 walpha0 = 1.033975766e-25 palpha0 = 7.395570986e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25 wub1 = 7.346839693e-40
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17 puc1 = 1.469367939e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.54 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.416818457e-01 lvth0 = -4.639353539e-8
+ k1 = 2.470831429e-01 lk1 = 9.210303897e-8
+ k2 = 6.961157274e-02 lk2 = -3.767169407e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.792280171e+04 lvsat = 2.104589919e-2
+ ua = -2.059561798e-09 lua = -4.034666577e-17
+ ub = 1.805365143e-18 lub = 1.010437038e-25
+ uc = 7.170268597e-11 luc = -7.785365576e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.204702371e-03 lu0 = 1.896620122e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.792502891e-01 lketa = -5.377655473e-08 wketa = 2.646977960e-23 pketa = -6.310887242e-30
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.980167143e+00 lags = 7.766315574e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.759934890e-01 lvoff = 1.677456896e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.037206100e+00 lnfactor = 8.280297364e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.361428571e-05 lcit = -3.547882857e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.918127253e-01 leta0 = 5.073405807e-08 weta0 = 3.308722450e-24 peta0 = -2.366582716e-30
+ etab = 2.237493824e-02 letab = -8.073894383e-9
+ dsub = 3.778380407e-01 ldsub = -7.421518127e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.417324086e+00 lpclm = -2.237365887e-07 ppclm = -1.009741959e-28
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 6.629674286e-03 lpdiblc2 = 1.481595881e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.984745545e-03 lalpha0 = -6.695024682e-10
+ alpha1 = 0.0
+ beta0 = 3.425952577e+01 lbeta0 = -1.127758428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.815118571e-01 lkt1 = -2.338054803e-8
+ kt2 = -3.436452571e-02 lkt2 = 2.574343801e-9
+ at = -3.756822857e+03 lat = 1.482731204e-2
+ ute = 9.931805714e-01 lute = -5.246609169e-7
+ ua1 = 4.886866343e-09 lua1 = -9.769024489e-16 pua1 = 1.880790961e-37
+ ub1 = -4.404562286e-18 lub1 = 9.239396537e-25
+ uc1 = -2.196574857e-12 luc1 = 2.455418768e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.55 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 2.473098676e-01 lvth0 = 9.713763628e-09 wvth0 = -1.657128471e-07 pvth0 = 3.158486865e-14
+ k1 = 1.274291442e+00 lk1 = -1.036828628e-07 wk1 = -1.603888740e-07 pk1 = 3.057011938e-14
+ k2 = -2.987896926e-01 lk2 = 3.254558710e-08 wk2 = 6.378621990e-08 pk2 = -1.215765351e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.439540464e+05 lvsat = 8.460343950e-03 wvsat = 8.962579389e-03 pvsat = -1.708267632e-9
+ ua = 8.570943735e-10 lua = -5.962613321e-16 wua = -3.898114521e-15 pua = 7.429806277e-22
+ ub = -1.705663686e-19 lub = 4.776562499e-25 wub = 2.470200726e-24 pub = -4.708202583e-31
+ uc = -8.480010875e-11 luc = 2.204406710e-17 wuc = 2.024523317e-16 puc = -3.858741443e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.205559967e-02 lu0 = -8.939160902e-09 wu0 = -6.435868652e-08 pu0 = 1.226676565e-14
+ a0 = 0.0
+ keta = 1.568280748e+00 lketa = -3.185257602e-07 wketa = -1.963466532e-06 pketa = 3.742367210e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.643310921e-01 lags = 1.582301938e-07 wags = 1.785819056e-08 pags = -3.403771121e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -3.404510258e-01 lvoff = 4.812017548e-08 wvoff = 3.410435352e-07 pvoff = -6.500289780e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.881776332e+00 lnfactor = -3.001283151e-07 wnfactor = -2.116930000e-06 pnfactor = 4.034868580e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.776689040e-01 leta0 = 4.803824572e-08 weta0 = 3.473644306e-07 peta0 = -6.620766046e-14
+ etab = -2.120138302e-01 letab = 3.660060488e-08 wetab = 1.304207654e-07 petab = -2.485819788e-14
+ dsub = 7.612804143e-01 ldsub = -8.050563453e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.828959136e+00 lpclm = -3.021942293e-07 wpclm = -1.812048274e-06 ppclm = 3.453764010e-13
+ pdiblc1 = 6.359752562e-01 lpdiblc1 = 6.938311616e-08 wpdiblc1 = 5.582865483e-07 ppdiblc1 = -1.064094161e-13
+ pdiblc2 = 7.268571389e-02 lpdiblc2 = -1.110868527e-08 wpdiblc2 = -1.903013432e-08 ppdiblc2 = 3.627143601e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.287806108e-04 lalpha0 = 6.544444824e-11 walpha0 = 1.658000174e-09 palpha0 = -3.160148331e-16
+ alpha1 = 0.0
+ beta0 = 2.253272867e+01 lbeta0 = 1.107369100e-06 wbeta0 = 1.202441081e-05 pbeta0 = -2.291852700e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 4.280353070e-01 lkt1 = -1.395602375e-07 wkt1 = -6.994830016e-07 pkt1 = 1.333214601e-13
+ kt2 = -4.304151645e-02 lkt2 = 4.228178236e-09 wkt2 = -4.157721604e-08 pkt2 = 7.924617378e-15
+ at = -9.260127561e+04 lat = 3.176106473e-02 wat = 1.484127250e-01 pat = -2.828746538e-8
+ ute = -2.207728711e+00 lute = 8.543239238e-08 wute = -1.015684588e-07 pute = 1.935894825e-14
+ ua1 = -4.255684850e-09 lua1 = 7.656678084e-16 wua1 = 2.946378216e-15 pua1 = -5.615796879e-22
+ ub1 = 6.546191676e-18 lub1 = -1.163274051e-24 wub1 = -5.070777404e-24 pub1 = 9.664901731e-31
+ uc1 = 4.677318984e-10 luc1 = -8.711294824e-17 wuc1 = -2.913117336e-16 puc1 = 5.552401642e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.56 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.57 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.58 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.058074269e-01 lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-01 pvsat = 4.235164736e-22
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16 puc = 4.701977403e-38
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.033923399e-01 lvoff = -2.743952297e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.365972934e+00 lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095731e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16 puc1 = -1.880790961e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.59 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.322046542e-01 lvth0 = 1.004565279e-8
+ k1 = 4.583847700e-01 lk1 = -9.143605620e-10
+ k2 = -2.429601160e-02 lk2 = -7.952904977e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.611812000e+02 lvsat = 8.411710788e-2
+ ua = -6.990916173e-10 lua = -8.205135605e-16
+ ub = 2.234268964e-18 lub = 9.853555799e-26
+ uc = 5.847047920e-11 luc = -1.408521648e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.438347102e-02 lu0 = -1.017317561e-8
+ a0 = 2.202768984e+00 la0 = -7.165335746e-7
+ keta = -2.506784320e-01 lketa = 1.396330174e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.136747526e+00 lags = 6.081310502e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.189493795e-01 lvoff = 3.839460957e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.867876868e-01 lnfactor = 1.613636150e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.672251120e-04 leta0 = -1.351628102e-10
+ etab = -5.283877540e-04 letab = 5.707641819e-11
+ dsub = 2.299473109e-01 ldsub = 3.464178733e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.573796660e-01 lpclm = -4.594153846e-08 wpclm = 2.117582368e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 8.771783000e-03 lpdiblc2 = 5.983981900e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.026313223e-04 lalpha0 = -1.572217669e-10
+ alpha1 = 0.0
+ beta0 = 2.161396292e+01 lbeta0 = -8.499367487e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.674992940e-01 lkt1 = -2.052231484e-9
+ kt2 = -5.161637500e-02 lkt2 = 2.920874017e-8
+ at = 1.947956140e+04 lat = 5.969961705e-2
+ ute = -1.146784080e+00 lute = 5.445525125e-8
+ ua1 = 2.097537420e-09 lua1 = -1.030179567e-16
+ ub1 = -2.064788220e-18 lub1 = 3.427836151e-25
+ uc1 = 3.200892914e-11 luc1 = -8.283476799e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.60 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.494846822e-01 lvth0 = -7.417543512e-9
+ k1 = 4.417433080e-01 lk1 = 1.590350094e-8
+ k2 = -2.483484439e-02 lk2 = -7.408360556e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.217170480e+04 lvsat = 1.175001425e-1
+ ua = -1.159636678e-09 lua = -3.550867226e-16
+ ub = 2.271786733e-18 lub = 6.062010003e-26
+ uc = 3.204681721e-11 luc = 1.261853632e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.758494212e-02 lu0 = -3.302582306e-9
+ a0 = 2.020313377e+00 la0 = -5.321439384e-7
+ keta = -2.274052120e-01 lketa = 1.161131012e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.282564612e+00 lags = -1.560431697e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.073091305e-01 lvoff = -7.924174767e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.187167452e+00 lnfactor = -1.047676407e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.891464901e-03 leta0 = 2.349589317e-09 weta0 = -4.135903063e-25 peta0 = -3.944304526e-31
+ etab = -8.261744920e-04 letab = 3.580196956e-10
+ dsub = 1.364052514e-01 ldsub = 4.409514786e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.659588400e-02 lpclm = 1.165465516e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.219616488e-02 lpdiblc2 = -7.582698428e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.870901370e-05 lalpha0 = 9.678277668e-11 palpha0 = 2.465190329e-32
+ alpha1 = 0.0
+ beta0 = 1.718699924e+01 lbeta0 = 3.623952740e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.683556200e-01 lkt1 = -1.186828428e-9
+ kt2 = -9.353640400e-03 lkt2 = -1.350197941e-8
+ at = 7.564972840e+04 lat = 2.934046279e-3
+ ute = -1.055830440e+00 lute = -3.746249734e-8
+ ua1 = 2.541635640e-09 lua1 = -5.518236178e-16
+ ub1 = -2.168290200e-18 lub1 = 4.473827161e-25
+ uc1 = -8.901892120e-11 luc1 = 3.947597756e-17 wuc1 = 4.930380658e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.61 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.092823266e-01 lvth0 = -3.795022070e-08 wvth0 = 4.235164736e-22
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.345075300e-01 lvoff = 5.963328048e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.817064934e+00 lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 6.203854594e-25 petab = -1.380506584e-30
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 palpha0 = 1.479114197e-31
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17 wuc1 = -1.232595164e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.62 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.416818457e-01 lvth0 = -4.639353539e-8
+ k1 = 2.470831429e-01 lk1 = 9.210303897e-8
+ k2 = 6.961157274e-02 lk2 = -3.767169407e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.792280171e+04 lvsat = 2.104589919e-2
+ ua = -2.059561798e-09 lua = -4.034666577e-17
+ ub = 1.805365143e-18 lub = 1.010437038e-25
+ uc = 7.170268597e-11 luc = -7.785365576e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.204702371e-03 lu0 = 1.896620122e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.792502891e-01 lketa = -5.377655473e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.980167143e+00 lags = 7.766315574e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.759934890e-01 lvoff = 1.677456896e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.037206100e+00 lnfactor = 8.280297364e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.361428571e-05 lcit = -3.547882857e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.918127253e-01 leta0 = 5.073405807e-08 weta0 = -1.323488980e-23 peta0 = 7.888609052e-30
+ etab = 2.237493824e-02 letab = -8.073894383e-09 petab = 3.155443621e-30
+ dsub = 3.778380407e-01 ldsub = -7.421518127e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.417324086e+00 lpclm = -2.237365887e-7
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 6.629674286e-03 lpdiblc2 = 1.481595881e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.984745545e-03 lalpha0 = -6.695024682e-10
+ alpha1 = 0.0
+ beta0 = 3.425952577e+01 lbeta0 = -1.127758428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.815118571e-01 lkt1 = -2.338054803e-8
+ kt2 = -3.436452571e-02 lkt2 = 2.574343801e-9
+ at = -3.756822857e+03 lat = 1.482731204e-2
+ ute = 9.931805714e-01 lute = -5.246609169e-7
+ ua1 = 4.886866343e-09 lua1 = -9.769024489e-16 pua1 = -3.761581923e-37
+ ub1 = -4.404562286e-18 lub1 = 9.239396537e-25 pub1 = -3.503246161e-46
+ uc1 = -2.196574857e-12 luc1 = 2.455418768e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.63 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -4.306389030e-01 lvth0 = 1.389307993e-07 wvth0 = 4.333565841e-07 pvth0 = -8.259776493e-14
+ k1 = 2.436557022e+00 lk1 = -3.252106824e-07 wk1 = -1.187424854e-06 pk1 = 2.263231772e-13
+ k2 = -2.287639682e-01 lk2 = 1.919868402e-08 wk2 = 1.907988488e-09 pk2 = -3.636626057e-16
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.269818083e+05 lvsat = 6.010071786e-02 wvsat = 2.483750474e-01 pvsat = -4.734028403e-8
+ ua = -1.087373226e-08 lua = 1.639634225e-15 wua = 6.467830437e-15 pua = -1.232768481e-21
+ ub = 3.109054962e-18 lub = -1.474395758e-25 wub = -4.278366632e-25 pub = 8.154566800e-32
+ uc = 2.809811888e-11 luc = 5.256649126e-19 wuc = 1.026898129e-16 puc = -1.957267834e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.777391381e-01 lu0 = 3.676571611e-08 wu0 = 1.475359335e-07 pu0 = -2.812034892e-14
+ a0 = 0.0
+ keta = -3.264023960e+00 lketa = 6.025115171e-07 wketa = 2.306599523e-06 pketa = -4.396378690e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.191679348e-01 lags = 1.668382916e-07 wags = 5.776661452e-08 pags = -1.101031673e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = 7.795543868e-01 lvoff = -1.653528562e-07 wvoff = -6.486492477e-07 pvoff = 1.236325466e-13
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.350922436e+01 lnfactor = -1.944519909e-06 wnfactor = -9.740574448e-06 pnfactor = 1.856553490e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.408013377e-01 leta0 = 6.007128758e-08 weta0 = 4.031514056e-07 peta0 = -7.684065790e-14
+ etab = 1.682800638e-01 letab = -3.588341132e-08 wetab = -2.056259341e-07 petab = 3.919230303e-14
+ dsub = 7.622193604e-01 ldsub = -8.068459766e-08 wdsub = -8.296997449e-10 pdsub = 1.581407714e-16
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.303974976e-01 lpclm = 9.031914504e-08 wpclm = 7.702215270e-09 ppclm = -1.468042230e-15
+ pdiblc1 = 2.478850522e+00 lpdiblc1 = -2.818689094e-07 wpdiblc1 = -1.070170180e-06 ppdiblc1 = 2.039744363e-13
+ pdiblc2 = 3.226476839e-01 lpdiblc2 = -5.875143675e-08 wpdiblc2 = -2.399090291e-07 ppdiblc2 = 4.572666095e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.308769144e-03 lalpha0 = 5.300414315e-10 walpha0 = 3.811941014e-09 palpha0 = -7.265559573e-16
+ alpha1 = 0.0
+ beta0 = -1.160575948e+02 lbeta0 = 2.752268474e-05 wbeta0 = 1.344897501e-04 pbeta0 = -2.563374637e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -9.494818413e-01 lkt1 = 1.229945309e-07 wkt1 = 5.177600265e-07 pkt1 = -9.868506104e-14
+ kt2 = -3.701330302e-01 lkt2 = 6.657182076e-08 wkt2 = 2.474572001e-07 pkt2 = -4.716534234e-14
+ at = 1.642598353e+05 lat = -1.719666302e-02 wat = -7.856259575e-02 pat = 1.497403075e-8
+ ute = -4.010255634e+00 lute = 4.289940238e-07 wute = 1.491234456e-06 pute = -2.842292874e-13
+ ua1 = -3.736743319e-09 lua1 = 6.667575527e-16 wua1 = 2.487815532e-15 pua1 = -4.741776404e-22
+ ub1 = 1.637036637e-19 lub1 = 5.322816369e-26 wub1 = 5.691081282e-25 pub1 = -1.084720092e-31
+ uc1 = 9.158292378e-10 luc1 = -1.725203011e-16 wuc1 = -6.872729475e-16 puc1 = 1.309942238e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.64 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.65 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.66 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.058074269e-01 lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-1
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.033923399e-01 lvoff = -2.743952297e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.365972934e+00 lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10 palpha0 = -4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095731e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.67 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.322046542e-01 lvth0 = 1.004565279e-8
+ k1 = 4.583847700e-01 lk1 = -9.143605620e-10
+ k2 = -2.429601160e-02 lk2 = -7.952904977e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.611812000e+02 lvsat = 8.411710788e-2
+ ua = -6.990916173e-10 lua = -8.205135605e-16
+ ub = 2.234268964e-18 lub = 9.853555799e-26
+ uc = 5.847047920e-11 luc = -1.408521648e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.438347102e-02 lu0 = -1.017317561e-08 wu0 = 1.323488980e-23
+ a0 = 2.202768984e+00 la0 = -7.165335746e-7
+ keta = -2.506784320e-01 lketa = 1.396330174e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.136747526e+00 lags = 6.081310502e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.189493795e-01 lvoff = 3.839460957e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.867876868e-01 lnfactor = 1.613636150e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.672251120e-04 leta0 = -1.351628102e-10
+ etab = -5.283877540e-04 letab = 5.707641819e-11
+ dsub = 2.299473109e-01 ldsub = 3.464178733e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.573796660e-01 lpclm = -4.594153846e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.771783000e-03 lpdiblc2 = 5.983981900e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.026313223e-04 lalpha0 = -1.572217669e-10
+ alpha1 = 0.0
+ beta0 = 2.161396292e+01 lbeta0 = -8.499367487e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.674992940e-01 lkt1 = -2.052231484e-9
+ kt2 = -5.161637500e-02 lkt2 = 2.920874017e-8
+ at = 1.947956140e+04 lat = 5.969961705e-2
+ ute = -1.146784080e+00 lute = 5.445525125e-8
+ ua1 = 2.097537420e-09 lua1 = -1.030179567e-16
+ ub1 = -2.064788220e-18 lub1 = 3.427836151e-25
+ uc1 = 3.200892914e-11 luc1 = -8.283476799e-17 puc1 = 5.877471754e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.68 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.494846822e-01 lvth0 = -7.417543512e-9
+ k1 = 4.417433080e-01 lk1 = 1.590350094e-8
+ k2 = -2.483484439e-02 lk2 = -7.408360556e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.217170480e+04 lvsat = 1.175001425e-1
+ ua = -1.159636678e-09 lua = -3.550867226e-16
+ ub = 2.271786733e-18 lub = 6.062010003e-26
+ uc = 3.204681721e-11 luc = 1.261853632e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.758494212e-02 lu0 = -3.302582306e-9
+ a0 = 2.020313377e+00 la0 = -5.321439384e-7
+ keta = -2.274052120e-01 lketa = 1.161131012e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.282564612e+00 lags = -1.560431697e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.073091305e-01 lvoff = -7.924174767e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.187167452e+00 lnfactor = -1.047676407e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.891464901e-03 leta0 = 2.349589317e-09 weta0 = 2.067951531e-25 peta0 = -2.958228395e-31
+ etab = -8.261744920e-04 letab = 3.580196956e-10
+ dsub = 1.364052514e-01 ldsub = 4.409514786e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.659588400e-02 lpclm = 1.165465516e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.219616488e-02 lpdiblc2 = -7.582698428e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.870901370e-05 lalpha0 = 9.678277668e-11 palpha0 = -1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.718699924e+01 lbeta0 = 3.623952740e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.683556200e-01 lkt1 = -1.186828428e-9
+ kt2 = -9.353640400e-03 lkt2 = -1.350197941e-8
+ at = 7.564972840e+04 lat = 2.934046279e-3
+ ute = -1.055830440e+00 lute = -3.746249734e-8
+ ua1 = 2.541635640e-09 lua1 = -5.518236178e-16
+ ub1 = -2.168290200e-18 lub1 = 4.473827161e-25
+ uc1 = -8.901892120e-11 luc1 = 3.947597756e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.69 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.092823266e-01 lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.345075300e-01 lvoff = 5.963328048e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.817064934e+00 lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 6.203854594e-25 petab = -5.176899691e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 palpha0 = 7.395570986e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.70 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.416818457e-01 lvth0 = -4.639353539e-8
+ k1 = 2.470831429e-01 lk1 = 9.210303897e-8
+ k2 = 6.961157274e-02 lk2 = -3.767169407e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.792280171e+04 lvsat = 2.104589919e-2
+ ua = -2.059561798e-09 lua = -4.034666577e-17
+ ub = 1.805365143e-18 lub = 1.010437038e-25
+ uc = 7.170268597e-11 luc = -7.785365576e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.204702371e-03 lu0 = 1.896620122e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.792502891e-01 lketa = -5.377655473e-08 pketa = -6.310887242e-30
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.980167143e+00 lags = 7.766315574e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.759934890e-01 lvoff = 1.677456896e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.037206100e+00 lnfactor = 8.280297364e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.361428571e-05 lcit = -3.547882857e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.918127253e-01 leta0 = 5.073405807e-08 weta0 = -9.926167351e-24 peta0 = 1.577721810e-30
+ etab = 2.237493824e-02 letab = -8.073894383e-09 petab = 1.577721810e-30
+ dsub = 3.778380407e-01 ldsub = -7.421518127e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.417324086e+00 lpclm = -2.237365887e-7
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 6.629674286e-03 lpdiblc2 = 1.481595881e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.984745545e-03 lalpha0 = -6.695024682e-10 walpha0 = -1.654361225e-24
+ alpha1 = 0.0
+ beta0 = 3.425952577e+01 lbeta0 = -1.127758428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.815118571e-01 lkt1 = -2.338054803e-8
+ kt2 = -3.436452571e-02 lkt2 = 2.574343801e-9
+ at = -3.756822857e+03 lat = 1.482731204e-2
+ ute = 9.931805714e-01 lute = -5.246609169e-7
+ ua1 = 4.886866343e-09 lua1 = -9.769024489e-16
+ ub1 = -4.404562286e-18 lub1 = 9.239396537e-25 wub1 = 7.346839693e-40 pub1 = -1.751623080e-46
+ uc1 = -2.196574857e-12 luc1 = 2.455418768e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.71 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 1.627290146e-01 lvth0 = 2.583487421e-08 wvth0 = 3.965890530e-09 pvth0 = -7.558987350e-16
+ k1 = 7.956742000e-01 lk1 = -1.245841652e-8
+ k2 = -2.177876132e-01 lk2 = 1.710659076e-08 wk2 = -6.035050807e-09 pk2 = 1.150280684e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.138888240e+05 lvsat = -4.869224657e-03 wvsat = 1.704014345e-03 pvsat = -3.247851342e-10
+ ua = -1.962922755e-09 lua = -5.876606748e-17 wua = 1.952313579e-17 pua = -3.721109681e-24
+ ub = 1.063189351e-19 lub = 4.248819110e-25 wub = 1.745093263e-24 pub = -3.326147759e-31
+ uc = 1.700034777e-10 luc = -2.652149647e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.685249332e-02 lu0 = -3.234488330e-10 wu0 = 6.719699428e-09 pu0 = -1.280774711e-15
+ a0 = 0.0
+ keta = 5.508284089e-01 lketa = -1.245993444e-07 wketa = -4.540183936e-07 pketa = 8.653590583e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.989946667e-01 lags = 1.516233165e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.168059176e-01 lvoff = 5.493417848e-09 wvoff = 1.886587311e-12 pvoff = -3.595835415e-19
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 7.137654675e-01 lnfactor = 4.942945556e-07 wnfactor = -4.811406220e-07 pnfactor = 9.170540255e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.163069406e-01 leta0 = -4.611355026e-08 weta0 = -1.058791184e-22
+ etab = -1.158710231e-01 letab = 1.827578585e-8
+ dsub = 7.610728120e-01 ldsub = -8.046606554e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.493419920e-01 lpclm = 1.320499657e-07 wpclm = 1.661413987e-07 ppclm = -3.166655059e-14
+ pdiblc1 = 1.0
+ pdiblc2 = -1.873215126e-02 lpdiblc2 = 6.315559830e-09 wpdiblc2 = 7.130488600e-09 ppdiblc2 = -1.359071127e-15
+ pdiblcb = 0.0
+ drout = -3.079223206e+01 ldrout = 6.535070191e-06 wdrout = 2.481166602e-05 pdrout = -4.729103544e-12
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.923300322e-03 lalpha0 = -4.671910087e-10 walpha0 = 2.575394538e-11 palpha0 = -4.908701990e-18
+ alpha1 = 0.0
+ beta0 = 6.162003200e+01 lbeta0 = -6.342670916e-06 wbeta0 = 5.913335496e-06 pbeta0 = -1.127081746e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.302269100e-01 lkt1 = 2.402454105e-08 wkt1 = 1.420011955e-07 pkt1 = -2.706542785e-14
+ kt2 = -2.817600667e-02 lkt2 = 1.394812071e-9
+ at = 1.193017444e+05 lat = -8.627650877e-03 wat = -4.602867321e-02 pat = 8.773065114e-9
+ ute = -1.949543333e+00 lute = 3.622225933e-8
+ ua1 = -2.988720667e-10 lua1 = 1.149929191e-17
+ ub1 = 9.501448000e-19 lub1 = -9.666751688e-26
+ uc1 = -3.390191333e-11 luc1 = 8.498456281e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.72 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.73 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 0.4215457
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.11023409
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.8262398
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.74 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.058074269e-01 lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-1
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-06 pags = 8.077935669e-28
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.033923399e-01 lvoff = -2.743952297e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.365972934e+00 lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10 palpha0 = -4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095730e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16 puc1 = -9.403954807e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.75 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.219859039e-01 lvth0 = 2.316514723e-07 wvth0 = 5.771604863e-08 pvth0 = -1.160438874e-13
+ k1 = 5.665343143e-01 lk1 = -2.183598343e-07 wk1 = -5.663250886e-08 pk1 = 1.138653223e-13
+ k2 = -7.557525680e-02 lk2 = 9.514914542e-08 wk2 = 2.685237675e-08 pk2 = -5.398938869e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.769825020e+04 lvsat = 1.005249695e-02 wvsat = -1.928973118e-02 pvsat = 3.878393351e-8
+ ua = 8.877692621e-10 lua = -4.011056045e-15 wua = -8.309596995e-16 pua = 1.670727572e-21
+ ub = 1.373510707e-19 lub = 4.314598673e-24 wub = 1.098051055e-24 pub = -2.207741450e-30
+ uc = -3.571360389e-11 luc = 1.752813010e-16 wuc = 4.931949511e-17 puc = -9.916177687e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.660410533e-02 lu0 = 5.468017040e-09 wu0 = 4.073664843e-09 pu0 = -8.190510533e-15
+ a0 = 2.524388491e+00 la0 = -1.363181755e-06 wa0 = -1.684160548e-07 pa0 = 3.386173198e-13
+ keta = -3.358443721e-01 lketa = 3.108676565e-07 wketa = 4.459714453e-08 pketa = -8.966701879e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.235109561e+00 lags = 4.103643429e-07 wags = -5.150727956e-08 pags = 1.035605363e-13
+ b0 = 2.717129478e-07 lb0 = -5.463060528e-13 wb0 = -1.422824851e-13 pb0 = 2.860731646e-19
+ b1 = 7.646430859e-08 lb1 = -1.537391389e-13 wb1 = -4.004053519e-14 pb1 = 8.050550006e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.920230222e-01 lvoff = 1.507613269e-07 wvoff = 3.826501297e-08 pvoff = -7.693563508e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.879069637e+00 lnfactor = 6.370428885e-06 wnfactor = 1.238881187e-06 pnfactor = -2.490894515e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.940003833e-05 lcit = -5.911171707e-11 wcit = -1.274932662e-11 pcit = 2.563379611e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.231202960e-03 leta0 = 3.480756672e-09 weta0 = 9.417468601e-10 peta0 = -1.893476237e-15
+ etab = 1.769534418e-03 letab = -4.563125901e-09 wetab = -1.203306945e-09 petab = 2.419368944e-15
+ dsub = -1.292870681e+00 ldsub = 3.408195727e-06 wdsub = 7.974236413e-07 pdsub = -1.603299973e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.149536981e-01 lpclm = -3.627598874e-07 wpclm = -8.251364191e-08 ppclm = 1.659019284e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -6.849276795e-03 lpdiblc2 = 3.739168472e-08 wpdiblc2 = 8.179967961e-09 ppdiblc2 = -1.644664358e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.039801412e-04 lalpha0 = -5.620537021e-10 walpha0 = -1.054363090e-10 palpha0 = 2.119902429e-16
+ alpha1 = 0.0
+ beta0 = 2.710697128e+01 lbeta0 = -1.189417936e-05 wbeta0 = -2.876413827e-06 pbeta0 = 5.783317641e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.993762807e-01 lkt1 = -1.390203619e-07 wkt1 = -3.567261589e-08 pkt1 = 7.172336151e-14
+ kt2 = -9.562608149e-02 lkt2 = 1.176946560e-07 wkt2 = 2.304568280e-08 pkt2 = -4.633564985e-14
+ at = 5.107714775e+04 lat = -3.830490064e-03 wat = -1.654607609e-02 pat = 3.326754059e-8
+ ute = -9.690507002e-01 lute = -3.028954822e-07 wute = -9.307008435e-08 pute = 1.871267116e-13
+ ua1 = 2.644858842e-09 lua1 = -1.203462407e-15 wua1 = -2.866048625e-16 pua1 = 5.762477365e-22
+ ub1 = -2.896969990e-18 lub1 = 2.015968282e-24 wub1 = 4.357719840e-25 pub1 = -8.761631510e-31
+ uc1 = 4.594796200e-10 luc1 = -9.423073390e-16 wuc1 = -2.238450273e-16 puc1 = 4.500628118e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.76 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 6.699221830e-01 lvth0 = -1.199729314e-07 wvth0 = -1.154320973e-07 pvth0 = 5.893962886e-14
+ k1 = 2.254442194e-01 lk1 = 1.263458156e-07 wk1 = 1.132650177e-07 pk1 = -5.783311805e-14
+ k2 = 7.772364600e-02 lk2 = -5.977472575e-08 wk2 = -5.370475349e-08 pk2 = 2.742164713e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.058458428e+05 lvsat = 1.551181573e-01 wvsat = 3.857946236e-02 pvsat = -1.969867348e-8
+ ua = -4.333358436e-09 lua = 1.265415607e-15 wua = 1.661919399e-15 pua = -8.485760451e-22
+ ub = 6.465622519e-18 lub = -2.080752452e-24 wub = -2.196102109e-24 pub = 1.121329737e-30
+ uc = 2.204149834e-10 luc = -8.356224933e-17 wuc = -9.863899022e-17 puc = 5.036506841e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.314367350e-02 lu0 = -1.124687055e-08 wu0 = -8.147329685e-09 pu0 = 4.160026537e-15
+ a0 = 1.377074363e+00 la0 = -2.037060979e-07 wa0 = 3.368321097e-07 pa0 = -1.719864752e-13
+ keta = -5.707333182e-02 lketa = 2.914164323e-08 wketa = -8.919428906e-08 pketa = 4.554260399e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.085840542e+00 lags = -1.459984387e-06 wags = 1.030145591e-07 pags = -5.259923388e-14
+ b0 = -5.434258956e-07 lb0 = 2.774732623e-13 wb0 = 2.845649702e-13 pb0 = -1.452988738e-19
+ b1 = -1.529286172e-07 lb1 = 7.808535193e-14 wb1 = 8.008107039e-14 pb1 = -4.088939454e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = 3.883815482e-02 lvoff = -8.254697863e-08 wvoff = -7.653002594e-08 pvoff = 3.907623125e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 6.918882099e+00 lnfactor = -2.520781139e-06 wnfactor = -2.477762375e-06 pnfactor = 1.265145469e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -4.369407667e-05 lcit = 2.486319555e-11 wcit = 2.549865325e-11 pcit = -1.301961235e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.705391244e-03 leta0 = 5.130345696e-10 weta0 = -1.883493720e-09 peta0 = 9.617118935e-16
+ etab = -5.422018836e-03 letab = 2.704657818e-09 wetab = 2.406613891e-09 petab = -1.228817053e-15
+ dsub = 3.182041234e+00 ldsub = -1.114150254e-06 wdsub = -1.594847283e-06 pdsub = 8.143290224e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.185521802e-01 lpclm = 2.774611532e-07 wpclm = 1.650272838e-07 ppclm = -8.426293111e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 5.343828447e-02 lpdiblc2 = -2.353492469e-08 wpdiblc2 = -1.635993592e-08 ppdiblc2 = 8.353383282e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.514066515e-04 lalpha0 = 3.024001905e-10 walpha0 = 2.108726180e-10 palpha0 = -1.076715588e-16
+ alpha1 = 0.0
+ beta0 = 6.200982523e+00 lbeta0 = 9.233412877e-06 wbeta0 = 5.752827655e-06 pbeta0 = -2.937393801e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.046016465e-01 lkt1 = 6.838039271e-08 wkt1 = 7.134523178e-08 pkt1 = -3.642887535e-14
+ kt2 = 7.866577258e-02 lkt2 = -5.844469168e-08 wkt2 = -4.609136561e-08 pkt2 = 2.353425128e-14
+ at = 1.245455570e+04 lat = 3.520150146e-02 wat = 3.309215218e-02 pat = -1.689685290e-8
+ ute = -1.411297200e+00 lute = 1.440388301e-07 wute = 1.861401687e-07 pute = -9.504317014e-14
+ ua1 = 1.446992797e-09 lua1 = 7.101018090e-18 wua1 = 5.732097250e-16 pua1 = -2.926808856e-22
+ ub1 = -5.039266595e-19 lub1 = -4.024413076e-25 wub1 = -8.715439680e-25 pub1 = 4.450103500e-31
+ uc1 = -9.439603029e-10 luc1 = 4.760090470e-16 wuc1 = 4.476900545e-16 puc1 = -2.285905418e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.77 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.092823266e-01 lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.345075300e-01 lvoff = 5.963328048e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.817064934e+00 lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 2.067951531e-25 petab = 4.437342592e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 palpha0 = 9.860761315e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-09 wkt2 = 2.646977960e-23
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.78 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 1.377874796e+00 lvth0 = -2.643054182e-07 wvth0 = -4.378724383e-07 pvth0 = 1.141095574e-13
+ k1 = -2.655009315e-01 lk1 = 2.256824487e-07 wk1 = 2.684146505e-07 pk1 = -6.994885793e-14
+ k2 = 3.237384768e-01 lk2 = -1.038971653e-07 wk2 = -1.330735533e-07 pk2 = 3.467896800e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.154821572e+05 lvsat = -1.480206885e-02 wvsat = -7.203295651e-02 pvsat = 1.877178847e-8
+ ua = 3.991792983e-09 lua = -1.617329722e-15 wua = -3.168791931e-15 pua = 8.257871773e-22
+ ub = -5.136743648e-19 lub = 7.053853995e-25 wub = 1.214365038e-24 pub = -3.164635289e-31
+ uc = -2.469399757e-10 luc = 7.525291205e-17 wuc = 1.668572298e-16 puc = -4.348299408e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.064451081e-01 lu0 = -2.448662961e-08 wu0 = -5.301453847e-08 pu0 = 1.381558872e-14
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.529171739e+00 lketa = -4.055660846e-07 wketa = -7.068863673e-07 pketa = 1.842145873e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.915880940e+00 lags = 7.598785728e-07 wags = -3.366347038e-08 pags = 8.772700380e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -6.259212383e-01 lvoff = 1.340257404e-07 wvoff = 2.356046659e-07 pvoff = -6.139857594e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -9.490229151e+00 lnfactor = 3.030887544e-06 wnfactor = 4.426425521e-06 pnfactor = -1.153526491e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 8.921245238e-05 lcit = -2.064276509e-11 wcit = -3.435047997e-11 pcit = 8.951735081e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.139505585e-01 leta0 = 5.650317738e-08 weta0 = 1.159247632e-08 peta0 = -3.020999329e-15
+ etab = -1.274041225e-01 letab = 3.095852884e-08 wetab = 7.843180514e-08 petab = -2.043932842e-14
+ dsub = 1.048788213e-01 ldsub = 6.371165444e-08 wdsub = 1.429350952e-07 pdsub = -3.724888581e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.305785655e+00 lpclm = -4.552696737e-07 wpclm = -4.652429008e-07 ppclm = 1.212422999e-13
+ pdiblc1 = -1.387891049e+01 lpdiblc1 = 3.718478074e-06 wpdiblc1 = 6.602162251e-06 ppdiblc1 = -1.720523483e-12
+ pdiblc2 = -2.039677038e-02 lpdiblc2 = 8.524687361e-09 wpdiblc2 = 1.415239775e-08 ppdiblc2 = -3.688114854e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.409091295e-03 lalpha0 = -7.800869707e-10 walpha0 = -2.222086520e-10 palpha0 = 5.790757471e-17
+ alpha1 = 0.0
+ beta0 = 3.758882952e+01 lbeta0 = -1.995374986e-06 wbeta0 = -1.743389910e-06 pbeta0 = 4.543274106e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 2.792496655e-01 lkt1 = -1.434550008e-07 wkt1 = -2.412777713e-07 pkt1 = 6.287698721e-14
+ kt2 = -1.537138301e-01 lkt2 = 3.367677254e-08 wkt2 = 6.249726327e-08 pkt2 = -1.628678681e-14
+ at = -6.024996399e+04 lat = 2.954942462e-02 wat = 2.958263335e-02 pat = -7.709234252e-9
+ ute = 1.226710045e+00 lute = -5.855186977e-07 wute = -1.222877087e-07 pute = 3.186817689e-14
+ ua1 = 6.937202640e-09 lua1 = -1.511220088e-15 wua1 = -1.073658602e-15 pua1 = 2.797954317e-22
+ ub1 = -7.751643142e-18 lub1 = 1.796188925e-24 wub1 = 1.752698890e-24 pub1 = -4.567533308e-31
+ uc1 = -2.179568168e-10 luc1 = 5.868253782e-17 wuc1 = 1.129828507e-16 puc1 = -2.944333089e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.79 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.644595440e+00 lvth0 = 3.117774088e-07 wvth0 = 9.503713413e-07 pvth0 = -1.504897070e-13
+ k1 = 1.991703707e+00 lk1 = -2.045407553e-07 wk1 = -6.263008512e-07 pk1 = 1.005839167e-13
+ k2 = -7.645738587e-01 lk2 = 1.035351659e-07 wk2 = 2.802895667e-07 pk2 = -4.410804268e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.561298815e+05 lvsat = -1.559695251e-01 wvsat = -3.869705154e-01 pvsat = 7.879888719e-8
+ ua = -1.474738778e-08 lua = 1.954358132e-15 wua = 6.714108247e-15 pua = -1.057893597e-21
+ ub = 2.238879825e-17 lub = -3.659825882e-24 wub = -9.923127033e-24 pub = 1.806342460e-30
+ uc = 1.522724601e-09 luc = -2.620451564e-16 wuc = -7.083524165e-16 puc = 1.233319645e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.521959802e-01 lu0 = 2.481036182e-08 wu0 = 9.524193260e-08 pu0 = -1.444209466e-14
+ a0 = 0.0
+ keta = -3.464776626e+00 lketa = 5.462804737e-07 wketa = 1.648753183e-06 pketa = -2.647703109e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.489935256e-01 lags = 1.757134998e-07 wags = 7.854809754e-08 pags = -1.261482447e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = 9.330548943e-01 lvoff = -1.631151105e-07 wvoff = -5.497577276e-07 pvoff = 8.829149626e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.228340739e+01 lnfactor = -1.119167582e-06 wnfactor = -6.539583617e-06 pnfactor = 9.365948509e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.748290556e-04 lcit = 2.968354632e-11 wcit = 8.015111994e-11 pcit = -1.287226986e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.679618846e-01 leta0 = -5.440933426e-08 weta0 = -2.704911141e-08 peta0 = 4.344087293e-15
+ etab = 2.336134519e-01 letab = -3.785142083e-08 wetab = -1.830075453e-07 petab = 2.939101178e-14
+ dsub = 1.397977657e+00 ldsub = -1.827529837e-07 wdsub = -3.335152222e-07 pdsub = 5.356254468e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.475975063e-01 lpclm = 1.457651569e-07 wpclm = 3.746878987e-07 ppclm = -3.884851045e-14
+ pdiblc1 = 3.041859114e+01 lpdiblc1 = -4.724625738e-06 wpdiblc1 = -1.540504525e-05 ppdiblc1 = 2.474050268e-12
+ pdiblc2 = -1.053046893e-01 lpdiblc2 = 2.470813671e-08 wpdiblc2 = 5.246419814e-08 ppdiblc2 = -1.099034401e-14
+ pdiblcb = 0.0
+ drout = 7.968756014e+01 ldrout = -1.452237820e-05 wdrout = -3.304107716e-05 pdrout = 6.297629308e-12
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.926154455e-03 lalpha0 = -3.068392089e-10 walpha0 = 5.479093787e-10 palpha0 = -8.887692195e-17
+ alpha1 = 0.0
+ beta0 = 3.798295661e+01 lbeta0 = -2.070495609e-06 wbeta0 = 1.829089003e-05 pbeta0 = -3.364206345e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -8.730433307e-01 lkt1 = 7.617204424e-08 wkt1 = 3.738820141e-07 pkt1 = -5.437246790e-14
+ kt2 = 2.503057037e-01 lkt2 = -4.332935061e-08 wkt2 = -1.458269476e-07 pkt2 = 2.341980779e-14
+ at = 2.383061371e+05 lat = -2.735536826e-02 wat = -1.083453235e-01 pat = 1.857983432e-8
+ ute = -2.494445438e+00 lute = 1.237335373e-07 wute = 2.853379870e-07 pute = -4.582528071e-14
+ ua1 = -7.896873311e-09 lua1 = 1.316154788e-15 wua1 = 3.978693352e-15 pua1 = -6.831828507e-22
+ ub1 = 8.760000131e-18 lub1 = -1.350930283e-24 wub1 = -4.089630744e-24 pub1 = 6.567946975e-31
+ uc1 = 4.695386512e-10 luc1 = -7.235409838e-17 wuc1 = -2.636266516e-16 puc1 = 4.233844025e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.80 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.263006254e-01 wvth0 = -2.061973410e-9
+ k1 = 6.583871577e-01 wk1 = -5.426139193e-8
+ k2 = -9.227296257e-02 wk2 = 1.505392322e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.548895758e+05 wvsat = -1.102943570e-1
+ ua = -4.970061183e-10 wua = -2.089443227e-16
+ ub = 2.678808214e-18 wub = -2.361389533e-25
+ uc = 1.571603771e-11 wuc = 2.877072299e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.428448092e-02 wu0 = -6.548236822e-9
+ a0 = 2.747888585e+00 wa0 = -3.607630987e-7
+ keta = 3.036500000e-01 wketa = -1.316778225e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.186027247e+00 wags = 1.197816429e-6
+ b0 = -1.303359231e-07 wb0 = 5.652017304e-14
+ b1 = -3.667858423e-08 wb1 = 1.590566805e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -6.369907348e-02 wvoff = -2.017990991e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.360202532e+00 wnfactor = -2.315529389e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.667117035e-01 weta0 = -8.096753024e-8
+ etab = -2.335038462e-01 wetab = 7.090344288e-8
+ dsub = 1.260730769e+00 wdsub = -3.038718981e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.657213846e-02 wpclm = 4.485149216e-8
+ pdiblc1 = 0.39
+ pdiblc2 = -1.577538731e-03 wpdiblc2 = 3.966439886e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.728345973e-05 walpha0 = 4.727582774e-11
+ alpha1 = 0.0
+ beta0 = 8.198856870e+00 wbeta0 = 4.160657583e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.625117577e-01 wkt1 = 2.116974223e-9
+ kt2 = -4.713656769e-02 wkt2 = 4.671523980e-9
+ at = -4.396644615e+03 wat = 2.715804444e-2
+ ute = -1.471369692e+00 wute = 1.260055471e-7
+ ua1 = 1.626314923e-09 wua1 = 1.462636736e-16
+ ub1 = -4.604513462e-19 wub1 = -4.360561737e-25
+ uc1 = 1.231856631e-10 wuc1 = -2.591824709e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.81 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.263006254e-01 wvth0 = -2.061973410e-9
+ k1 = 6.583871577e-01 wk1 = -5.426139193e-8
+ k2 = -9.227296257e-02 wk2 = 1.505392322e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.548895758e+05 wvsat = -1.102943570e-1
+ ua = -4.970061183e-10 wua = -2.089443227e-16
+ ub = 2.678808214e-18 wub = -2.361389533e-25
+ uc = 1.571603771e-11 wuc = 2.877072299e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.428448092e-02 wu0 = -6.548236822e-9
+ a0 = 2.747888585e+00 wa0 = -3.607630987e-7
+ keta = 3.036500000e-01 wketa = -1.316778225e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.186027247e+00 wags = 1.197816429e-6
+ b0 = -1.303359231e-07 wb0 = 5.652017304e-14
+ b1 = -3.667858423e-08 wb1 = 1.590566805e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -6.369907348e-02 wvoff = -2.017990991e-8
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.360202532e+00 wnfactor = -2.315529389e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.667117035e-01 weta0 = -8.096753024e-8
+ etab = -2.335038462e-01 wetab = 7.090344288e-8
+ dsub = 1.260730769e+00 wdsub = -3.038718981e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.657213846e-02 wpclm = 4.485149216e-8
+ pdiblc1 = 0.39
+ pdiblc2 = -1.577538731e-03 wpdiblc2 = 3.966439886e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.728345972e-05 walpha0 = 4.727582774e-11
+ alpha1 = 0.0
+ beta0 = 8.198856870e+00 wbeta0 = 4.160657583e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.625117577e-01 wkt1 = 2.116974223e-9
+ kt2 = -4.713656769e-02 wkt2 = 4.671523980e-9
+ at = -4.396644615e+03 wat = 2.715804444e-2
+ ute = -1.471369692e+00 wute = 1.260055471e-7
+ ua1 = 1.626314923e-09 wua1 = 1.462636736e-16
+ ub1 = -4.604513462e-19 wub1 = -4.360561737e-25
+ uc1 = 1.231856631e-10 wuc1 = -2.591824709e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.82 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.738013783e-01 lvth0 = 2.105534805e-07 wvth0 = 1.387942298e-08 pvth0 = -6.393456435e-14
+ k1 = 9.110024564e-01 lk1 = -1.013138917e-06 wk1 = -1.309680274e-07 pk1 = 3.076396321e-13
+ k2 = -1.905525136e-01 lk2 = 3.941599674e-07 wk2 = 4.489650890e-08 pk2 = -1.196866741e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.842381770e+05 lvsat = -2.123005500e+00 wvsat = -2.710310598e-01 pvsat = 6.446506201e-7
+ ua = -6.658331792e-11 lua = -1.726253683e-15 wua = -3.396422060e-16 pua = 5.241769308e-22
+ ub = 2.179121203e-18 lub = 2.004044727e-24 wub = -8.440899235e-26 pub = -6.085281813e-31
+ uc = -8.191765585e-11 luc = 3.915696914e-16 wuc = 3.252354335e-17 puc = -1.189001368e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.381667481e-02 lu0 = 1.876183179e-09 wu0 = -6.406187497e-09 pu0 = -5.697030224e-16
+ a0 = 2.981205791e+00 la0 = -9.357419897e-07 wa0 = -4.316098686e-07 pa0 = 2.841380552e-13
+ keta = 9.113955274e-01 lketa = -2.437424212e-06 wketa = -3.162197519e-07 pketa = 7.401238621e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -5.080268189e+00 lags = 1.160764272e-05 wags = 2.076652690e-06 pags = -3.524660712e-12
+ b0 = -1.303359231e-07 wb0 = 5.652017304e-14
+ b1 = -3.667858423e-08 wb1 = 1.590566805e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -4.087657400e-02 lvoff = -9.153191642e-08 wvoff = -2.710996188e-08 pvoff = 2.779366642e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.160627715e+00 lnfactor = -7.220785238e-06 wnfactor = -7.782520456e-07 pnfactor = 2.192591437e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.333108837e-01 leta0 = -1.069222672e-06 weta0 = -1.619203713e-07 peta0 = 3.246694644e-13
+ etab = -4.665685383e-01 letab = 9.347292543e-07 wetab = 1.416735367e-07 petab = -2.838305381e-13
+ dsub = 1.789760525e+00 ldsub = -2.121726737e-06 wdsub = -4.645117833e-07 pdsub = 6.442623235e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.922244887e-02 lpclm = 4.644057719e-07 wpclm = 8.001251860e-08 ppclm = -1.410168127e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -1.559126595e-02 lpdiblc2 = 5.620345440e-08 wpdiblc2 = 8.221708157e-09 ppdiblc2 = -1.706617893e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.446134850e-04 lalpha0 = 1.112259799e-09 walpha0 = 1.314870899e-10 palpha0 = -3.377376880e-16
+ alpha1 = 0.0
+ beta0 = -3.195732937e+00 lbeta0 = 4.569914188e-05 wbeta0 = 7.620624778e-06 pbeta0 = -1.387654443e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.259927002e-01 lkt1 = -1.464633321e-07 wkt1 = -8.972037591e-09 pkt1 = 4.447359078e-14
+ kt2 = -4.470531731e-02 lkt2 = -9.750772796e-09 wkt2 = 3.933274800e-09 pkt2 = 2.960822160e-15
+ at = 2.597889468e+04 lat = -1.218241379e-01 wat = 1.793451193e-02 pat = 3.699189948e-8
+ ute = -1.676265414e+00 lute = 8.217547833e-07 wute = 1.882221331e-07 pute = -2.495258399e-13
+ ua1 = 1.348984707e-09 lua1 = 1.112260566e-15 wua1 = 2.304749938e-16 pua1 = -3.377379208e-22
+ ub1 = 9.758307782e-19 lub1 = -5.760353088e-24 wub1 = -8.721832408e-25 pub1 = 1.749131215e-30
+ uc1 = 3.666732095e-10 luc1 = -9.765311535e-16 wuc1 = -9.985324055e-17 puc1 = 2.965236848e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.83 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.381617257e-01 lvth0 = -1.199094340e-07 wvth0 = -3.602859651e-08 pvth0 = 3.641049964e-14
+ k1 = 3.337479079e-01 lk1 = 1.474890783e-07 wk1 = 4.431531627e-08 pk1 = -4.478505862e-14
+ k2 = 5.418406536e-02 lk2 = -9.790739830e-08 wk2 = -2.941775331e-08 pk2 = 2.972958149e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.367288279e+05 lvsat = 3.318707601e-01 wvsat = 9.971557125e-02 pvsat = -1.007725563e-7
+ ua = -6.624486809e-10 lua = -5.282067842e-16 wua = -1.587076885e-16 pua = 1.603899900e-22
+ ub = 4.464093734e-18 lub = -2.590121044e-24 wub = -7.782409013e-25 pub = 7.864902549e-31
+ uc = 2.014080279e-10 luc = -1.780849284e-16 wuc = -5.350830054e-17 puc = 5.407548852e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.701376392e-02 lu0 = -4.476388418e-08 wu0 = -1.344998360e-08 pu0 = 1.359255343e-14
+ a0 = 3.481936494e+00 la0 = -1.942511141e-06 wa0 = -5.836567466e-07 pa0 = 5.898435081e-13
+ keta = -4.735943648e-01 lketa = 3.472364651e-07 wketa = 1.043324289e-07 pketa = -1.054383526e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.840867191e-01 lags = 2.165500258e-06 wags = 6.506571873e-07 pags = -6.575541535e-13
+ b0 = -3.184448869e-07 lb0 = 3.782118827e-13 wb0 = 1.136394599e-13 pb0 = -1.148440382e-19
+ b1 = -8.961541325e-08 lb1 = 1.064347884e-13 wb1 = 3.197993618e-14 pb1 = -3.231892351e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -4.218182329e-02 lvoff = -8.890758221e-08 wvoff = -2.671362293e-08 pvoff = 2.699678734e-14
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -4.699993891e-01 lnfactor = 2.089553618e-06 wnfactor = 6.278378746e-07 pnfactor = -6.344929560e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.987362739e-03 leta0 = -2.954200816e-09 weta0 = -8.876341556e-10 peta0 = 8.970430777e-16
+ etab = -3.353448808e-03 letab = 3.388995365e-09 wetab = 1.018274730e-09 petab = -1.029068443e-15
+ dsub = 1.214009774e+00 ldsub = -9.641222777e-07 wdsub = -2.896850679e-07 pdsub = 2.927557296e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.788877482e-01 lpclm = 6.608540962e-08 wpclm = 1.985635724e-08 ppclm = -2.006683463e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 1.324891407e-02 lpdiblc2 = -1.782611562e-09 wpdiblc2 = -5.356125082e-10 ppdiblc2 = 5.412900008e-16
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.300344155e-04 lalpha0 = -2.441872695e-10 walpha0 = -7.336974508e-11 palpha0 = 7.414746438e-17
+ alpha1 = 0.0
+ beta0 = 1.714064457e+01 lbeta0 = 4.810821258e-06 wbeta0 = 1.445483747e-06 pbeta0 = -1.460805875e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.425955310e-01 lkt1 = 8.797831968e-08 wkt1 = 2.643441200e-08 pkt1 = -2.671461677e-14
+ kt2 = -6.754671257e-02 lkt2 = 3.617413653e-08 wkt2 = 1.086906447e-08 pkt2 = -1.098427656e-14
+ at = -1.555344175e+05 lat = 2.431265275e-01 wat = 7.305102916e-02 pat = -7.382537007e-8
+ ute = -1.480946619e+00 lute = 4.290468132e-07 wute = 1.289135809e-07 pute = -1.302800648e-13
+ ua1 = 1.694184417e-09 lua1 = 4.182020280e-16 wua1 = 1.256551017e-16 pua1 = -1.269870458e-22
+ ub1 = -1.881744825e-18 lub1 = -1.491157961e-26 wub1 = -4.480408814e-27 pub1 = 4.527901147e-33
+ uc1 = -2.775289966e-10 luc1 = 3.187018019e-16 wuc1 = 9.575875931e-17 puc1 = -9.677380216e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.84 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 4.037349415e-01 lvth0 = 1.594227410e-8
+ k1 = 4.866341600e-01 lk1 = -7.017768096e-9
+ k2 = -4.611989947e-02 lk2 = 3.459788568e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.688132680e+04 lvsat = 1.096928755e-1
+ ua = -5.009604218e-10 lua = -6.914068188e-16
+ ub = 1.401395356e-18 lub = 5.050419372e-25
+ uc = -7.047233185e-12 luc = 3.257995846e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.435587300e-02 lu0 = -1.653819614e-9
+ a0 = 2.153811616e+00 la0 = -6.003081391e-7
+ keta = -2.627560000e-01 lketa = 1.341632136e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.323392852e+00 lags = -1.581278596e-6
+ b0 = 1.127829600e-07 lb0 = -5.758697938e-14
+ b1 = 3.173890360e-08 lb1 = -1.620588418e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.376406321e-01 lvoff = 7.563089958e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.205144350e+00 lnfactor = 3.966533552e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.510600000e-05 lcit = -5.160123600e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.637958740e-03 leta0 = 2.730749071e-09 weta0 = -1.550963649e-25 peta0 = -1.232595164e-32
+ etab = 1.276500000e-04 letab = -1.290030900e-10
+ dsub = -4.956880000e-01 ldsub = 7.636982928e-07 pdsub = -5.048709793e-29
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.620019160e-01 lpclm = 8.315023169e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.571215528e-02 lpdiblc2 = -4.271963126e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.486711313e-05 lalpha0 = 5.410880632e-11
+ alpha1 = 0.0
+ beta0 = 1.946704422e+01 lbeta0 = 2.459761774e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.400790320e-01 lkt1 = -1.562485426e-8
+ kt2 = -2.762124600e-02 lkt2 = -4.174539992e-9
+ at = 8.876529520e+04 lat = -3.762762129e-3
+ ute = -9.820566400e-01 lute = -7.513139962e-8
+ ua1 = 2.768818520e-09 lua1 = -6.678231963e-16
+ ub1 = -2.513713280e-18 lub1 = 6.237557408e-25
+ uc1 = 8.841616320e-11 luc1 = -5.112237653e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.85 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 5.092823266e-01 lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.345075300e-01 lvoff = 5.963328048e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 1.817064934e+00 lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = -6.203854594e-25 petab = 1.602373714e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 walpha0 = -5.169878828e-26 palpha0 = -2.465190329e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17 puc1 = -7.346839693e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.86 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 3.681378229e-01 lvth0 = -1.167963037e-9
+ k1 = 3.534651714e-01 lk1 = 6.437988233e-8
+ k2 = 1.686991157e-02 lk2 = -2.392721717e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.937364457e+04 lvsat = 2.848580954e-2
+ ua = -3.315463863e-09 lua = 2.869414123e-16
+ ub = 2.286660094e-18 lub = -2.438176057e-26
+ uc = 1.378339890e-10 luc = -2.501918314e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.580679657e-02 lu0 = 7.372216747e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = -1.009132772e-01 lketa = 1.923407063e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.993509143e+00 lags = 7.801084826e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -8.261519446e-02 lvoff = -7.559814600e-9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 7.171397426e-01 lnfactor = 3.708472098e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.872182252e-01 leta0 = 4.953673133e-08 weta0 = -8.271806126e-24 peta0 = -2.761013168e-30
+ etab = 5.346018086e-02 letab = -1.617470861e-08 petab = 7.888609052e-31
+ dsub = 4.344881727e-01 ldsub = -2.218454253e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.232932200e+00 lpclm = -1.756840633e-7
+ pdiblc1 = 1.345722857e+00 lpdiblc1 = -2.490613766e-7
+ pdiblc2 = 1.223876000e-02 lpdiblc2 = 1.986814400e-11
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.896676555e-03 lalpha0 = -6.465516894e-10
+ alpha1 = 0.0
+ beta0 = 3.356855993e+01 lbeta0 = -9.476927294e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.771386000e-01 lkt1 = 1.539781160e-9
+ kt2 = -9.594694286e-03 lkt2 = -3.880674269e-9
+ at = 7.967800000e+03 lat = 1.177187532e-2
+ ute = 9.447137143e-01 lute = -5.120304539e-7
+ ua1 = 4.461338229e-09 lua1 = -8.660098224e-16 wua1 = -7.888609052e-31
+ ub1 = -3.709906971e-18 lub1 = 7.429124788e-25 wub1 = -3.673419846e-40
+ uc1 = 4.258244457e-11 luc1 = -9.213993695e-18 wuc1 = -3.081487911e-33
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.87 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.363696e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 2.666245949e-01 lvth0 = 1.818045821e-08 wvth0 = 1.215707731e-07 pvth0 = -2.317138935e-14
+ k1 = 5.474494667e-01 lk1 = 2.740647565e-8
+ k2 = -1.908607291e-01 lk2 = 1.566624293e-08 wk2 = 3.149886801e-08 pk2 = -6.003684242e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.527559666e+04 lvsat = 4.652595492e-02 wvsat = 4.728897020e-02 pvsat = -9.013277720e-9
+ ua = 7.879959843e-11 lua = -3.600052035e-16 wua = 2.847320897e-16 pua = -5.426993629e-23
+ ub = -4.769423026e-18 lub = 1.320507682e-24 wub = 1.854035626e-24 pub = -3.533791902e-31
+ uc = -4.060716821e-10 luc = 7.864923778e-17 wuc = 1.280700919e-16 puc = -2.441015952e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.740901945e-02 lu0 = -6.582717787e-09 wu0 = 4.346724492e-09 pu0 = -8.284856881e-16
+ a0 = 0.0
+ keta = -5.173987401e-01 lketa = 9.861619987e-08 wketa = 3.706227627e-07 pketa = -7.064069856e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.301260000e-01 lags = 1.466236244e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre)
+ voff = -3.347005338e-01 lvoff = 4.048765109e-08 wvoff = 4.413854116e-12 pvoff = -8.412805944e-19
*(mismatch parameter sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -4.591715034e+00 lnfactor = 1.382714930e-06 wnfactor = 7.783132240e-07 pnfactor = -1.483465005e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.055864403e-01 leta0 = -4.439183791e-8
+ etab = -1.884032559e-01 letab = 2.992446244e-8
+ dsub = 6.288891707e-01 ldsub = -5.923737274e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.643546667e-02 lpclm = 5.618021405e-8
+ pdiblc1 = -5.105553333e+00 lpdiblc1 = 9.805518653e-07 wpdiblc1 = 2.646977960e-22 ppdiblc1 = -8.835242138e-29
+ pdiblc2 = 1.567812667e-02 lpdiblc2 = -6.356751427e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.740867895e-03 lalpha0 = -8.074545589e-10 walpha0 = -6.726911048e-10 palpha0 = 1.282149246e-16
+ alpha1 = 0.0
+ beta0 = 1.723718178e+02 lbeta0 = -2.740359367e-05 wbeta0 = -3.998683961e-05 pbeta0 = 7.621491630e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.086873333e-02 lkt1 = -4.921125543e-8
+ kt2 = -8.597228000e-02 lkt2 = 1.067689357e-8
+ at = -1.419322429e+05 lat = 4.034282350e-02 wat = 5.654505002e-02 pat = -1.077748653e-8
+ ute = -1.836454000e+00 lute = 1.806011240e-8
+ ua1 = 2.642099863e-09 lua1 = -5.192629900e-16 wua1 = -5.915323654e-16 pua1 = 1.127460689e-22
+ ub1 = -6.707176000e-19 lub1 = 1.636429846e-25
+ uc1 = -1.383862920e-10 luc1 = 2.527864750e-17 wuc1 = 6.162975822e-33 puc1 = -1.469367939e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -0.3015
+ k1 = 0.64774
+ k2 = 0.002296
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.00225441
+ a0 = 1.75737
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.283503
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -0.3015
+ k1 = 0.64774
+ k2 = 0.002296
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.00225441
+ a0 = 1.75737
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.283503
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.058359263e-01 lvth0 = 3.451288897e-8
+ k1 = 0.64774
+ k2 = -9.370912500e-05 lk2 = 1.902148721e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.063707319e-09 lua = 4.641116804e-16
+ ub = 3.130202425e-18 lub = -7.028652274e-25
+ uc = 3.789249356e-11 luc = 9.122276612e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.176779101e-03 lu0 = 6.179225463e-10
+ a0 = 1.849196603e+00 la0 = -7.309167992e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.705724364e-01 lags = 1.029240538e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 9.025288750e-05 lpdiblc2 = 1.398008393e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.927296312e-03 ldelta = 6.131159568e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112493750e-01 lkt1 = 7.879655016e-8
+ kt2 = -0.055045
+ at = 2.990532506e+05 lat = -1.070845117e-1
+ ute = -3.115370919e-01 lute = 7.070414446e-7
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.751307275e-19 lub1 = 2.108595682e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.628429926e-01 lvth0 = -1.357283800e-7
+ k1 = 0.64774
+ k2 = -1.128156000e-02 lk2 = 6.332257971e-08 pk2 = 2.524354897e-29
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.561076335e+05 lvsat = -1.280885418e-1
+ ua = -3.110237112e-09 lua = 6.483580312e-16
+ ub = 3.171996025e-18 lub = -8.683574350e-25
+ uc = 4.861983037e-11 luc = 4.874519417e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.036878354e-03 lu0 = 1.171894531e-9
+ a0 = 2.218745970e+00 la0 = -2.194239909e-6
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.422712694e-01 lags = -1.809854002e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.221488000e-04 lpdiblc2 = 1.306183409e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.970993700e-02 ldelta = 6.735784214e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.761903100e+05 lat = -4.125279825e-1
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.565136819e-19 lub1 = 1.371407218e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.398697895e-01 lvth0 = 1.522488522e-8
+ k1 = 0.64774
+ k2 = 1.089799375e-01 lk2 = -1.723598900e-7
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 90748.0
+ ua = -2.247467100e-09 lua = -1.042455501e-15
+ ub = 1.852758050e-18 lub = 1.717019187e-24
+ uc = 7.920646150e-11 luc = -1.119695617e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.930255010e-03 lu0 = -5.789003708e-10
+ a0 = 9.687460835e-01 la0 = 2.554473696e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.459449270e-01 lags = 2.037651493e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.040698600e-03 lpdiblc2 = 1.965217428e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.711239350e-02 ldelta = 1.182632009e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 2.048988850e+05 lat = -7.683961238e-2
+ ute = -0.13298
+ ua1 = 7.976886000e-10 lua1 = -1.991078563e-16
+ ub1 = -3.072346025e-19 lub1 = 4.325160460e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.094349710e-01 lvth0 = -2.920234108e-8
+ k1 = 0.64774
+ k2 = -4.248662200e-02 lk2 = 4.874342021e-08 pk2 = -2.524354897e-29
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.005122150e+04 lvsat = 1.017122415e-3
+ ua = -3.146447850e-09 lua = 2.698316490e-16
+ ub = 3.137067850e-18 lub = -1.577520440e-25
+ uc = 5.217208400e-11 luc = 2.826647638e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.824002460e-03 lu0 = 1.035951789e-9
+ a0 = 1.056633090e+00 la0 = 1.271543119e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -2.318686300e-02 lags = 4.506552798e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -1.539712750e-01 lvoff = -4.076895632e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.595652800e+00 lnfactor = -8.518049980e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 9.396700000e-04 lpdiblc2 = 1.384183122e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.075824550e-02 ldelta = 2.110178763e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.489350000e-01 lkt1 = 8.405970375e-8
+ kt2 = -9.202608700e-02 lkt2 = 5.398314175e-8
+ at = 2.025317050e+05 lat = -7.338412137e-2
+ ute = 4.956445000e-02 lute = -2.664692609e-7
+ ua1 = 6.6129e-10
+ ub1 = -1.051962950e-20 lub1 = -6.136358374e-28
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.362382505e-01 lvth0 = -3.477893583e-9
+ k1 = 0.64774
+ k2 = 2.549013300e-02 lk2 = -1.649727040e-08 wk2 = -2.646977960e-23 pk2 = -6.310887242e-30
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.467314300e+04 lvsat = -3.418766744e-3
+ ua = -2.795142150e-09 lua = -6.733399654e-17
+ ub = 2.835418650e-18 lub = 1.317557757e-25
+ uc = 9.281615400e-11 luc = -1.074166980e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.917118940e-03 lu0 = -1.316675266e-11
+ a0 = 1.274688670e+00 la0 = -8.212453103e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.698134110e-01 lags = -2.250173321e-8
+ b0 = 7.194076050e-08 lb0 = -6.904514489e-14
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -2.098287250e-01 lvoff = 1.284023132e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.478947200e+00 lnfactor = 2.682769980e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.007644950e-02 lpdiblc2 = 3.401205191e-08 ppdiblc2 = -1.262177448e-29
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.216615250e-02 ldelta = 1.015304889e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -4.964241050e-01 lkt1 = -6.231262773e-8
+ kt2 = -1.717199800e-02 lkt2 = -1.785807017e-8
+ at = 1.874319130e+05 lat = -5.889209600e-2
+ ute = -7.139720000e-02 lute = -1.503763173e-7
+ ua1 = 4.451523300e-10 lua1 = 2.074381288e-16
+ ub1 = 5.295630895e-19 lub1 = -5.189580254e-25 wub1 = 4.591774808e-41 pub1 = 3.503246161e-46
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.620328200e-01 lvth0 = 8.381159745e-9
+ k1 = 0.64774
+ k2 = -3.375434500e-02 lk2 = 1.074037836e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.428050850e+04 lvsat = -3.238253033e-3
+ ua = -3.060750500e-09 lua = 5.477944238e-17
+ ub = 3.039400000e-18 lub = 3.797535000e-26
+ uc = 8.249041000e-11 luc = -5.994408998e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.319304050e-03 lu0 = 2.616786430e-10
+ a0 = 1.294423900e+00 la0 = -9.119780303e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.120937500e-01 lags = 4.034880938e-9
+ b0 = -2.398025350e-07 lb0 = 7.427883522e-14
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.416210500e-02 lpdiblc2 = 5.887793202e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.684411500e-02 ldelta = 8.002355629e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.526100000e-01 lkt1 = 9.493837500e-9
+ kt2 = -0.056015
+ at = 1.297958650e+05 lat = -3.239392293e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.178348025e-01 wvth0 = 1.151505243e-7
+ k1 = 0.64774
+ k2 = 2.535185090e-04 wk2 = 1.439826494e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.123303443e-09 wua = 8.311482974e-16
+ ub = 3.234534534e-18 wub = -1.357957497e-24
+ uc = 5.089054169e-11 wuc = -1.083874332e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.277990689e-03 wu0 = -1.662296595e-10
+ a0 = 1.762570880e+00 wa0 = -3.666307265e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.111731961e-01 wags = -1.950582250e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.357346608e-03 wpdiblc2 = -3.600456115e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.354475070e-03 wdelta = 7.243626489e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.178348025e-01 wvth0 = 1.151505243e-7
+ k1 = 0.64774
+ k2 = 2.535185090e-04 wk2 = 1.439826494e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.123303443e-09 wua = 8.311482974e-16
+ ub = 3.234534534e-18 wub = -1.357957497e-24
+ uc = 5.089054169e-11 wuc = -1.083874332e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.277990689e-03 wu0 = -1.662296595e-10
+ a0 = 1.762570880e+00 wa0 = -3.666307265e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.111731961e-01 wags = -1.950582250e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.357346608e-03 wpdiblc2 = -3.600456115e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.354475070e-03 wdelta = 7.243626489e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.900797910e-01 lvth0 = -2.209229527e-07 wvth0 = -1.110712680e-07 pvth0 = 1.800668911e-12
+ k1 = 0.64774
+ k2 = 1.834052690e-02 lk2 = -1.439680650e-07 wk2 = -1.299502666e-07 pk2 = 1.148978224e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.328819191e-09 lua = 1.635853976e-15 wua = 1.868879105e-15 pua = -8.260077794e-21
+ ub = 3.545774003e-18 lub = -2.477388364e-24 wub = -2.929529449e-24 pub = 1.250931985e-29
+ uc = 1.049570611e-11 luc = 3.215327925e-16 wuc = 1.931308587e-16 puc = -1.623547039e-21
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.017186517e-03 lu0 = 2.075936007e-09 wu0 = 1.125031646e-09 pu0 = -1.027811717e-14
+ a0 = 2.092105355e+00 la0 = -2.623012041e-06 wa0 = -1.712360477e-06 pa0 = 1.333813241e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.540913612e-01 lags = -3.416178644e-07 wags = -5.887581414e-07 pags = 3.133752910e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.080502740e-04 lpdiblc2 = 1.962394283e-08 wpdiblc2 = 1.397917910e-09 ppdiblc2 = -3.978580764e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.202606045e-02 ldelta = 1.224252176e-07 wdelta = 1.265603573e-07 pdelta = -4.308142442e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112493750e-01 lkt1 = 7.879655016e-8
+ kt2 = -0.055045
+ at = 2.990532506e+05 lat = -1.070845117e-1
+ ute = -3.115370919e-01 lute = 7.070414446e-7
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.751307275e-19 lub1 = 2.108595682e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.473509370e-01 lvth0 = -7.860935325e-07 wvth0 = -8.141494660e-07 pvth0 = 4.584682806e-12
+ k1 = 0.64774
+ k2 = -7.395726696e-02 lk2 = 2.215081242e-07 wk2 = 4.418260033e-07 pk2 = -1.115112861e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.377756714e+05 lvsat = -4.514735550e-01 wvsat = -5.757105034e-01 pvsat = 2.279669666e-6
+ ua = -3.639276963e-09 lua = 2.865189138e-15 wua = 3.729412466e-15 pua = -1.562732477e-20
+ ub = 3.986487150e-18 lub = -4.222502247e-24 wub = -5.741672105e-24 pub = 2.364470173e-29
+ uc = 6.639541898e-11 luc = 1.001839045e-16 wuc = -1.253071987e-16 puc = -3.626119416e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.284907704e-03 lu0 = 4.975577035e-09 wu0 = 5.300940392e-09 pu0 = -2.681367183e-14
+ a0 = 3.424311646e+00 la0 = -7.898215898e-06 wa0 = -8.498512260e-06 pa0 = 4.020959693e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.892182002e-01 lags = -8.766863652e-07 wags = -1.035887400e-06 pags = 4.904272991e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.444947878e-03 lpdiblc2 = 9.514708398e-09 wpdiblc2 = -1.496445557e-08 ppdiblc2 = 2.500510075e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.338684151e-02 ldelta = -5.739852094e-08 wdelta = -9.641394332e-08 pdelta = 4.521082425e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 5.786534212e+05 lat = -1.214231287e+00 wat = -1.427243051e+00 pat = 5.651525671e-6
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -2.439533039e-19 lub1 = 4.833797650e-25 wub1 = 6.163966964e-25 pub1 = -2.440776819e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -8.952321824e-01 lvth0 = 6.795667381e-07 wvth0 = 3.914970542e-06 pvth0 = -4.683210129e-12
+ k1 = 0.64774
+ k2 = 2.815367481e-01 lk2 = -4.751712719e-07 wk2 = -1.216421636e-06 pk2 = 2.134637950e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.845648890e+05 lvsat = 7.681583582e-01 wvsat = 3.350669729e+00 pvsat = -5.415053994e-6
+ ua = -5.072658005e-10 lua = -3.272769738e-15 wua = -1.226737156e-14 pua = 1.572237272e-20
+ ub = -7.882126803e-19 lub = 5.134715744e-24 wub = 1.861725378e-23 pub = -2.409270328e-29
+ uc = 2.333871217e-10 luc = -2.270780849e-16 wuc = -1.086880838e-15 puc = 1.521831997e-21
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 6.095460906e-03 lu0 = -4.451904602e-09 wu0 = -2.231279611e-08 pu0 = 2.730234828e-14
+ a0 = -1.379631464e+00 la0 = 1.516311611e-06 wa0 = 1.655464799e-05 pa0 = -8.888333860e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.500989599e-01 lags = -1.191972434e-06 wags = -3.553982431e-06 pags = 9.839109728e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -6.473021715e-03 lpdiblc2 = 2.699169931e-08 wpdiblc2 = 2.419581170e-08 ppdiblc2 = -5.173923304e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.447425998e-03 ldelta = 2.066668481e-08 wdelta = 1.660825445e-07 pdelta = -6.231924940e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.124757619e-01 lkt1 = 4.333512119e-07 wkt1 = 1.558803504e-06 pkt1 = -3.054865167e-12
+ kt2 = -2.051672798e-01 lkt2 = 2.942021378e-07 wkt2 = 1.058271699e-06 pkt2 = -2.073947962e-12
+ at = -8.405999133e+05 lat = 1.567150435e+00 wat = 7.370137138e+00 pat = -1.158914015e-5
+ ute = -0.13298
+ ua1 = 8.435353413e-10 lua1 = -2.889560076e-16 wua1 = -3.231919265e-16 pua1 = 6.333753779e-22
+ ub1 = 4.252388548e-20 lub1 = -7.804390684e-26 wub1 = -2.465586786e-24 pub1 = 3.599140310e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -4.951140259e-01 lvth0 = 9.549425915e-08 wvth0 = 1.308925558e-06 pvth0 = -8.790359643e-13
+ k1 = 0.64774
+ k2 = -1.828955162e-01 lk2 = 2.027837260e-07 wk2 = 9.897981781e-07 pk2 = -1.085891424e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.190611777e+05 lvsat = -4.049347925e-01 wvsat = -2.319322127e+00 pvsat = 2.861716617e-6
+ ua = -3.206959457e-09 lua = 6.681080769e-16 wua = 4.265704008e-16 pua = -2.807609054e-21
+ ub = 3.110224872e-18 lub = -5.560284719e-25 wub = 1.892268388e-25 pub = 2.807609054e-30
+ uc = 4.266515319e-11 luc = 5.132830861e-17 wuc = 6.701813906e-17 puc = -1.625720340e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.775068428e-03 lu0 = 1.854788317e-09 wu0 = 3.449554645e-10 pu0 = -5.772304582e-15
+ a0 = -1.497635286e+00 la0 = 1.688567689e-06 wa0 = 1.800605438e-05 pa0 = -1.100702434e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.423560121e+00 lags = 1.835051409e-06 wags = 9.871788445e-06 pags = -9.759159307e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -8.345965092e-02 lvoff = -1.436982996e-07 wvoff = -4.970645018e-07 pvoff = 7.255899064e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.742976056e+00 lnfactor = -3.002356225e-07 wnfactor = -1.038540265e-06 pnfactor = 1.516009152e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.741299014e-02 lpdiblc2 = -7.875906499e-09 wpdiblc2 = -1.161269901e-07 ppdiblc2 = 1.530969768e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.520137611e-03 ldelta = 3.197033833e-09 wdelta = 3.692550728e-08 pdelta = 1.262177356e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.216556273e-01 lkt1 = 1.548015204e-07 wkt1 = -1.923031553e-07 pkt1 = -4.986872209e-13
+ kt2 = 5.809619276e-02 lkt2 = -9.009671626e-08 wkt2 = -1.058271699e-06 pkt2 = 1.015676263e-12
+ at = 9.217763381e+05 lat = -1.005478298e+00 wat = -5.070241678e+00 pat = 6.570702823e-6
+ ute = 3.300117136e-01 lute = -6.758521539e-07 wute = -1.976984379e-06 pute = 2.885902947e-12
+ ua1 = 5.192954496e-10 lua1 = 1.843531742e-16 wua1 = 1.000976099e-15 pua1 = -1.299578898e-21
+ ub1 = -9.458320519e-21 lub1 = -2.162881622e-27 wub1 = -7.481589408e-27 pub1 = 1.092125014e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.436049725e-01 lvth0 = -4.991655480e-08 wvth0 = 5.193095541e-08 pvth0 = 3.273646055e-13
+ k1 = 0.64774
+ k2 = 5.859115358e-02 lk2 = -2.898310533e-08 wk2 = -2.333422682e-07 pk2 = 8.801761978e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.729136042e+04 lvsat = -7.692121042e-02 wvsat = 1.225311034e-01 pvsat = 5.181479794e-7
+ ua = -1.814808597e-09 lua = -6.680087105e-16 wua = -6.910761385e-15 pua = 4.234395127e-21
+ ub = 1.545566720e-18 lub = 9.456521889e-25 wub = 9.092679615e-24 pub = -5.737479748e-30
+ uc = 9.889274851e-11 luc = -2.636125998e-18 wuc = -4.283633319e-17 puc = -5.713920428e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 4.490833180e-03 lu0 = -7.516669036e-10 wu0 = -1.109373802e-08 pu0 = 5.205981487e-15
+ a0 = 1.049581319e+00 la0 = -7.561234469e-07 wa0 = 1.586871311e-06 pa0 = 4.751286610e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.647098407e-01 lags = 1.187593136e-07 wags = 7.409168983e-07 pags = -9.958053407e-13
+ b0 = 1.276335481e-06 lb0 = -1.224962978e-12 wb0 = -8.490257731e-12 pb0 = 8.148524858e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -2.803403491e-01 lvoff = 4.525795049e-08 wvoff = 4.970645018e-07 pvoff = -2.285254047e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.331623944e+00 lnfactor = 9.455956666e-08 wnfactor = 1.038540265e-06 pnfactor = -4.774688868e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.820576011e-02 lpdiblc2 = 4.550418905e-08 wpdiblc2 = 1.278007260e-07 ppdiblc2 = -8.101264862e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.231590859e-03 ldelta = 4.433716578e-09 wdelta = 1.264278630e-07 pdelta = 4.031784975e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.172493476e-01 lkt1 = -1.373524065e-07 wkt1 = -1.263074176e-06 pkt1 = 5.289852666e-13
+ kt2 = -1.717199800e-02 lkt2 = -1.785807017e-8
+ at = -2.961663665e+05 lat = 1.634422130e-01 wat = 3.409076744e+00 pat = -1.567323033e-6
+ ute = -3.518444636e-01 lute = -2.144068786e-08 wute = 1.976984379e-06 pute = -9.089185683e-13
+ ua1 = 5.413001391e-10 lua1 = 1.632341736e-16 wua1 = -6.777841728e-16 pua1 = 3.116112735e-22
+ ub1 = 5.285017805e-19 lub1 = -5.184700886e-25 wub1 = 7.481589408e-27 pub1 = -3.439660730e-33
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -5.351597619e-01 lvth0 = 3.815075964e-08 wvth0 = 1.220440718e-06 pvth0 = -2.098577580e-13
+ k1 = 0.64774
+ k2 = 2.265497763e-03 lk2 = -3.087385067e-09 wk2 = -2.539182075e-07 pk2 = 9.747740787e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.859804205e+05 lvsat = 1.820429908e-01 wvsat = 4.090490232e+00 pvsat = -1.306121230e-6
+ ua = -4.060526255e-09 lua = 3.644599824e-16 wua = 7.047817205e-15 pua = -2.183061379e-21
+ ub = 4.511979923e-18 lub = -4.181562813e-25 wub = -1.038080197e-23 pub = 3.215453409e-30
+ uc = 1.551521309e-10 luc = -2.850137704e-17 wuc = -5.122213897e-16 puc = 1.586605755e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.117949080e-03 lu0 = 3.392665616e-10 wu0 = 1.419431325e-09 pu0 = -5.469481180e-16
+ a0 = -3.888856237e+00 la0 = 1.514323219e-06 wa0 = 3.653900463e-05 pa0 = -1.131795668e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.054057549e+00 lags = -1.981682952e-07 wags = -4.525458319e-06 pags = 1.425410665e-12
+ b0 = -4.254451602e-06 lb0 = 1.317816384e-12 wb0 = 2.830085910e-11 pb0 = -8.766191108e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.364520468e-01 lpdiblc2 = 9.067291935e-08 wpdiblc2 = 4.391065910e-07 ppdiblc2 = -2.241355201e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.407641743e-03 ldelta = 5.272277184e-09 wdelta = 1.722624257e-07 pdelta = 1.924540953e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.037045606e-01 lkt1 = -5.654622351e-09 wkt1 = -3.447539066e-07 pkt1 = 1.067875226e-13
+ kt2 = -0.056015
+ at = 1.297958650e+05 lat = -3.239392293e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.933528311e-01 wvth0 = -8.468693289e-9
+ k1 = 0.64774
+ k2 = 1.012318950e-02 wk2 = -3.543763201e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.111169900e-09 wua = 7.698812081e-16
+ ub = 3.072328930e-18 wub = -5.389168457e-25
+ uc = 3.016401799e-11 wuc = 9.381772402e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.905656756e-03 wu0 = 1.713832557e-9
+ a0 = 1.759731627e+00 wa0 = -2.232655504e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.900699199e-01 wags = -8.849938464e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.244490933e-04 wpdiblc2 = 4.644693329e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.317621807e-02 wdelta = 2.284237544e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 2.899606391e+05 wat = -2.201860255e-2
+ ute = -1.174447810e-01 wute = -5.315259861e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.463681985e-19 wub1 = -1.147123000e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.933528311e-01 wvth0 = -8.468693289e-9
+ k1 = 0.64774
+ k2 = 1.012318950e-02 wk2 = -3.543763201e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.111169900e-09 wua = 7.698812081e-16
+ ub = 3.072328930e-18 wub = -5.389168457e-25
+ uc = 3.016401799e-11 wuc = 9.381772402e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.905656756e-03 wu0 = 1.713832557e-9
+ a0 = 1.759731627e+00 wa0 = -2.232655504e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.900699199e-01 wags = -8.849938464e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.244490933e-04 wpdiblc2 = 4.644693329e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.317621807e-02 wdelta = 2.284237544e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 2.899606391e+05 wat = -2.201860255e-2
+ ute = -1.174447810e-01 wute = -5.315259861e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.463681985e-19 wub1 = -1.147123000e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.958342625e-01 lvth0 = 1.975157389e-08 wvth0 = -8.201465116e-08 pvth0 = 5.854074382e-13
+ k1 = 0.64774
+ k2 = -9.778015386e-04 lk2 = 8.836111340e-08 wk2 = -3.240433758e-08 pk2 = -2.414426533e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.156450601e-09 lua = 3.604230637e-16 wua = 9.985214917e-16 pua = -1.819919497e-21
+ ub = 3.072328930e-18 wub = -5.389168457e-25
+ uc = 3.016401799e-11 wuc = 9.381772402e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.723062933e-03 lu0 = 1.453401181e-09 wu0 = 2.610178682e-09 pu0 = -7.134691068e-15
+ a0 = 1.839346741e+00 la0 = -6.337164009e-07 wa0 = -4.360816335e-07 pa0 = 3.293386986e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.364234381e-01 lags = 4.270125842e-07 wags = 5.394034202e-09 pags = -7.473681406e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.513579764e-03 lpdiblc2 = 1.781415019e-08 wpdiblc2 = 8.494995703e-09 ppdiblc2 = -3.064744433e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.180500002e-02 ldelta = 1.091455284e-08 wdelta = 6.227848174e-09 pdelta = 1.322474834e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112493750e-01 lkt1 = 7.879655016e-8
+ kt2 = -0.055045
+ at = 3.077306500e+05 lat = -1.414448437e-01 wat = -4.381564292e-02 pat = 1.734989920e-7
+ ute = -1.020658852e-01 lute = -1.224121660e-07 wute = -1.057703492e-06 pute = 4.188241402e-12
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.706099845e-19 lub1 = 1.929585561e-25 wub1 = -2.282703075e-26 pub1 = 9.038933501e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.562254245e-01 lvth0 = 2.588854773e-07 wvth0 = 2.405409533e-07 pvth0 = -6.918321165e-13
+ k1 = 0.64774
+ k2 = 1.761123283e-02 lk2 = 1.475318454e-08 wk2 = -2.053979644e-08 pk2 = -7.112488210e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.918974676e-09 lua = -5.799222339e-16 wua = 9.231953519e-17 pua = 1.768413700e-21
+ ub = 2.778925643e-18 lub = 1.161803665e-24 wub = 3.557865500e-25 pub = -3.542801771e-30
+ uc = -2.490208249e-12 luc = 1.293025723e-16 wuc = 2.225237496e-16 puc = -5.096436848e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.270770451e-03 lu0 = -7.153836651e-10 wu0 = 3.229270096e-10 pu0 = 1.922253743e-15
+ a0 = 1.334565902e+00 la0 = 1.365089524e-06 wa0 = 2.053445716e-06 pa0 = -6.564518938e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.780976250e-01 lags = 2.619932225e-07 wags = 3.014441000e-08 pags = -8.453734412e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.408670462e-03 lpdiblc2 = 1.739873559e-08 wpdiblc2 = 4.493997166e-09 ppdiblc2 = -1.480449037e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.266166368e-02 ldelta = 7.522378933e-09 wdelta = 8.235728198e-09 pdelta = 1.242967805e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 2.848968128e+05 lat = -5.102855685e-02 wat = 5.605098002e-02 pat = -2.219478681e-7
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.678553806e-02 lvth0 = -4.063318401e-07 wvth0 = -5.206561873e-07 pvth0 = 7.999239797e-13
+ k1 = 0.64774
+ k2 = 5.025413836e-02 lk2 = -4.921874958e-08 wk2 = -4.858368854e-08 pk2 = -1.616586457e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.157275256e+05 lvsat = -7.681583582e-01 wvsat = -1.195264989e+00 pvsat = 2.342420561e-6
+ ua = -3.009981238e-09 lua = -4.015721230e-16 wua = 3.698347649e-16 pua = 1.224553229e-21
+ ub = 2.903708702e-18 lub = 9.172600652e-25 wub = -2.472665970e-26 pub = -2.797091008e-30
+ uc = -3.224380557e-11 luc = 1.876121847e-16 wuc = 2.543954352e-16 puc = -5.721042207e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 9.146796540e-04 lu0 = 1.942215275e-09 wu0 = 3.847030380e-09 pu0 = -4.984107836e-15
+ a0 = 2.005699166e+00 la0 = 4.983611068e-08 wa0 = -5.392337249e-07 pa0 = -1.483515403e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -3.616324866e-01 lags = 1.515704309e-06 wags = 1.554652311e-06 pags = -3.833027801e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.195305916e-03 lpdiblc2 = 2.873909442e-08 wpdiblc2 = 2.784291210e-08 ppdiblc2 = -6.056252642e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.454495035e-02 ldelta = 6.084054077e-08 wdelta = 2.069701677e-07 pdelta = -2.651730373e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.702242381e-01 lkt1 = -4.333512119e-07 wkt1 = -6.743004561e-07 pkt1 = 1.321460319e-12
+ kt2 = 9.507727976e-02 lkt2 = -2.942021378e-07 wkt2 = -4.577825797e-07 pkt2 = 8.971394105e-13
+ at = 1.100532716e+06 lat = -1.649471019e+00 wat = -2.431414080e+00 pat = 4.652861783e-6
+ ute = -0.13298
+ ua1 = 9.067491425e-10 lua1 = -4.128392545e-16 wua1 = -6.423835679e-16 pua1 = 1.258911197e-21
+ ub1 = -9.396030676e-19 lub1 = 1.602532782e-24 wub1 = 2.493563087e-24 pub1 = -4.886760259e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.400441623e-01 lvth0 = -8.043006338e-08 wvth0 = 2.097629888e-08 pvth0 = 9.275958033e-15
+ k1 = 0.64774
+ k2 = 1.178609028e-01 lk2 = -1.479077240e-07 wk2 = -5.288406828e-07 pk2 = 6.848892828e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.903544755e+05 lvsat = 4.085198429e-01 wvsat = 1.262799853e+00 pvsat = -1.245739592e-6
+ ua = -3.166649539e-09 lua = -1.728755708e-16 wua = 2.230295818e-16 pua = 1.438852095e-21
+ ub = 3.637729034e-18 lub = -1.542261147e-25 wub = -2.474351625e-24 pub = 7.787490349e-31
+ uc = 1.880736170e-10 luc = -1.339961729e-16 wuc = -6.672070671e-16 puc = 7.732050320e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.010540999e-03 lu0 = -1.117218323e-09 wu0 = -5.893437261e-09 pu0 = 9.234539802e-15
+ a0 = 2.394186849e+00 la0 = -5.172587843e-07 wa0 = -1.645304523e-06 pa0 = 1.310714442e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 9.797326015e-01 lags = -4.423533787e-07 wags = -2.263393022e-06 pags = 1.740363875e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 6.714228767e+00 lnfactor = -6.097271768e-06 wnfactor = -2.109097576e-05 pnfactor = 3.078755187e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.406441466e-02 lpdiblc2 = 3.876627591e-08 wpdiblc2 = 4.281495479e-08 ppdiblc2 = -8.241796572e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.790876938e-02 ldelta = -1.572877660e-08 wdelta = -1.266175852e-07 pdelta = 2.217816850e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.518139565e-01 lkt1 = 2.696493796e-07 wkt1 = 9.698578519e-07 pkt1 = -1.078599771e-12
+ kt2 = -2.421483668e-01 lkt2 = 1.980629998e-07 wkt2 = 4.577825797e-07 pkt2 = -4.393568308e-13
+ at = -6.358975664e+05 lat = 8.852830864e-01 wat = 2.795073820e+00 pat = -2.976503929e-6
+ ute = -6.632089890e-01 lute = 7.740017667e-07 wute = 3.038182250e-06 pute = -4.434986540e-12
+ ua1 = 5.903123375e-10 lua1 = 4.907937160e-17 wua1 = 6.423835679e-16 pua1 = -6.165276293e-22
+ ub1 = 4.828937376e-19 lub1 = -4.739569296e-25 wub1 = -2.493563087e-24 pub1 = 2.393197173e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.275042699e-01 lvth0 = 3.509774930e-09 wvth0 = -2.936790011e-08 pvth0 = 5.759380302e-14
+ k1 = 0.64774
+ k2 = -5.698295111e-02 lk2 = 1.989866482e-08 wk2 = 3.502373848e-07 pk2 = -1.588058926e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.909500921e+04 lvsat = 9.233069989e-02 wvsat = 3.153996828e-01 pvsat = -3.364722780e-7
+ ua = -3.837572347e-09 lua = 4.710425946e-16 wua = 3.302977849e-15 pua = -1.517128254e-21
+ ub = 3.978470502e-18 lub = -4.812527382e-25 wub = -3.192019875e-24 pub = 1.467531137e-30
+ uc = 4.437997240e-11 luc = 3.913802512e-18 wuc = 2.324203695e-16 puc = -9.021240019e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 7.616481119e-04 lu0 = 1.041156625e-09 wu0 = 7.736401608e-09 pu0 = -3.846698053e-15
+ a0 = 1.689496340e+00 la0 = 1.590679314e-07 wa0 = -1.644314317e-06 pa0 = 1.301210942e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.335959417e-01 lags = -1.101487195e-07 wags = -6.167960424e-07 pags = 1.600424235e-13
+ b0 = -1.318902119e-06 lb0 = 1.265816309e-12 wb0 = 4.614129815e-12 pb0 = -4.428411089e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 3.612495872e-01 wnfactor = 1.098774460e-5
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.163536690e-03 lpdiblc2 = 3.214315827e-08 wpdiblc2 = -2.894381490e-08 ppdiblc2 = -1.354748652e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.747194670e-03 ldelta = 1.705779472e-08 wdelta = 1.288737721e-07 pdelta = -2.342614519e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.368988850e-01 lkt1 = -3.259036032e-08 wkt1 = -1.539762416e-07 pkt1 = -1.615587134e-27
+ kt2 = -1.010471396e-02 lkt2 = -2.464089603e-08 wkt2 = -3.568552991e-08 pkt2 = 3.424918733e-14
+ at = 5.003923223e+05 lat = -2.052711343e-01 wat = -6.130651057e-01 pat = 2.944574051e-7
+ ute = 5.911019272e-01 lute = -4.298231351e-07 wute = -2.784327241e-06 pute = 1.153166944e-12
+ ua1 = 4.070694500e-10 lua1 = 2.249467329e-16
+ ub1 = 4.795829717e-19 lub1 = -4.707794221e-25 wub1 = 2.544921246e-25 pub1 = -2.442488166e-31
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.985272472e-01 lvth0 = -5.578741128e-08 wvth0 = -4.793508287e-07 pvth0 = 2.644734544e-13
+ k1 = 0.64774
+ k2 = -3.423243876e-03 lk2 = -4.725410586e-09 wk2 = -2.251934869e-07 pk2 = 1.057484507e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.335596538e+05 lvsat = -1.809744204e-01 wvsat = -1.562513180e+00 pvsat = 5.268981605e-7
+ ua = -2.881034865e-09 lua = 3.127448699e-17 wua = 1.092095741e-15 pua = -5.006752053e-22
+ ub = 2.752719524e-18 lub = 8.228627404e-26 wub = -1.497596022e-24 pub = 6.885197713e-31
+ uc = -8.003748206e-12 luc = 2.799721806e-17 wuc = 3.116175797e-16 puc = -1.266233176e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.523871802e-03 lu0 = 6.907242834e-10 wu0 = 4.419163943e-09 pu0 = -2.321598036e-15
+ a0 = 5.729119855e+00 la0 = -1.698148980e-06 wa0 = -1.202598461e-05 pa0 = 4.903094012e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -6.795654428e-02 lags = 2.123900360e-07 wags = 1.140037398e-06 pags = -6.476617509e-13
+ b0 = 4.396340397e-06 lb0 = -1.361766438e-12 wb0 = -1.538043272e-11 pb0 = 4.764089033e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 3.612495872e-01 wnfactor = 1.098774460e-5
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.097044619e-02 lpdiblc2 = 3.849088492e-08 wpdiblc2 = -1.440059720e-07 ppdiblc2 = 3.935234022e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.786927005e-02 ldelta = -7.824829430e-09 wdelta = -1.077854093e-07 pdelta = 8.537791347e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.729718544e-01 lkt1 = 2.996918734e-08 wkt1 = 5.004227853e-09 pkt1 = -7.309127084e-14
+ kt2 = -7.957261347e-02 lkt2 = 7.296970774e-09 wkt2 = 1.189517664e-07 pkt2 = -3.684530963e-14
+ at = 1.131592643e+05 lat = -2.724073588e-02 wat = 8.400481814e-02 pat = -2.602049242e-8
+ ute = -2.308989607e-01 lute = -5.190822693e-08 wute = -8.461833648e-07 pute = 2.621052972e-13
+ ua1 = 8.9635e-10
+ ub1 = -4.312183725e-19 lub1 = -5.203850413e-26 wub1 = -8.483070821e-25 pub1 = 2.627631187e-31
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.114931867e-01 wvth0 = 4.684847086e-8
+ k1 = 0.64774
+ k2 = -1.062828730e-02 wk2 = 2.784187983e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.844218308e-09 wua = -4.416044384e-17
+ ub = 2.872303364e-18 wub = 7.104071401e-26
+ uc = 5.901170046e-11 wuc = 5.849658793e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.489161177e-03 wu0 = -6.550465836e-11
+ a0 = 1.872875643e+00 wa0 = -3.673476921e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.448266893e-01 wags = -2.554745677e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.696427525e-03 wpdiblc2 = -1.368653756e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.473866424e-02 wdelta = -1.241612479e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.908560200e-01 wkt1 = -3.200032162e-8
+ kt2 = -0.055045
+ at = 2.871894475e+05 wat = -1.356813637e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.114931867e-01 wvth0 = 4.684847086e-8
+ k1 = 0.64774
+ k2 = -1.062828730e-02 wk2 = 2.784187983e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.844218308e-09 wua = -4.416044384e-17
+ ub = 2.872303364e-18 wub = 7.104071401e-26
+ uc = 5.901170046e-11 wuc = 5.849658793e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.489161177e-03 wu0 = -6.550465836e-11
+ a0 = 1.872875643e+00 wa0 = -3.673476921e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.448266893e-01 wags = -2.554745677e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.696427525e-03 wpdiblc2 = -1.368653756e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.473866424e-02 wdelta = -1.241612479e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.908560200e-01 wkt1 = -3.200032162e-8
+ kt2 = -0.055045
+ at = 2.871894475e+05 wat = -1.356813637e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.489798341e-01 lvth0 = 2.983843416e-07 wvth0 = 8.004734853e-08 pvth0 = -2.642547665e-13
+ k1 = 0.64774
+ k2 = -2.910344165e-02 lk2 = 1.470576098e-07 wk2 = 5.336193312e-08 pk2 = -2.031332442e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.824908567e-09 lua = -1.537007083e-16 wua = -1.248212545e-17 pua = -2.521514948e-22
+ ub = 2.915415159e-18 lub = -3.431591099e-25 wub = -6.042430730e-26 pub = 1.046428703e-30
+ uc = 5.901170046e-11 wuc = 5.849658793e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.667052143e-03 lu0 = -1.415967615e-09 wu0 = -2.684201268e-10 pu0 = 1.615156400e-15
+ a0 = 1.832789622e+00 la0 = 3.190747085e-07 wa0 = -4.160863688e-07 pa0 = 3.879476823e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.384334850e-01 lags = 5.088830839e-08 wags = -3.056751988e-07 pags = 3.995844738e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.864751278e-03 lpdiblc2 = -1.339814998e-09 wpdiblc2 = -4.856278219e-09 ppdiblc2 = 2.776061882e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.940244608e-02 ldelta = 4.247496246e-08 wdelta = -1.693978866e-08 pdelta = 3.600723346e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.903670107e-01 lkt1 = -3.892391985e-09 wkt1 = -6.367864001e-08 pkt1 = 2.521514948e-13
+ kt2 = -0.055045
+ at = 3.022161518e+05 lat = -1.196088098e-01 wat = -2.699974336e-02 pat = 1.069122338e-7
+ ute = -4.489223769e-01 lute = 1.251052827e-6
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.521398367e-19 lub1 = 1.599779781e-26 wub1 = -7.914986241e-26 pub1 = 6.300131173e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.901567753e-01 lvth0 = 6.545973451e-08 wvth0 = 3.907134669e-08 pvth0 = -1.020000433e-13
+ k1 = 0.64774
+ k2 = 9.356532334e-03 lk2 = -5.234272139e-09 wk2 = 4.632070755e-09 pk2 = -1.017517169e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.838017356e-09 lua = -1.017931809e-16 wua = -1.545515533e-16 pua = 3.104079223e-22
+ ub = 2.797647912e-18 lub = 1.231697489e-25 wub = 2.986949021e-25 pub = -3.755935860e-31
+ uc = 7.357684716e-11 luc = -5.767433966e-17 wuc = -9.434977028e-18 puc = 6.052333669e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.390057084e-03 lu0 = -3.191364314e-10 wu0 = -4.082541032e-11 pu0 = 7.139382213e-16
+ a0 = 2.161300974e+00 la0 = -9.817481187e-07 wa0 = -4.675985585e-07 pa0 = 5.919230752e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.010784530e-01 lags = -1.971701038e-07 wags = -3.448730810e-07 pags = 5.547982877e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 5.084365503e-05 lpdiblc2 = 9.802555713e-09 wpdiblc2 = 4.335773577e-11 ppdiblc2 = 8.359285348e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.225946006e-02 ldelta = 7.075940138e-08 wdelta = 9.462207101e-09 pdelta = -6.853806924e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.032778113e+05 lat = -1.238127156e-1
+ ute = -1.439208871e-01 lute = 4.332317780e-08 wute = 3.336311932e-08 pute = -1.321096117e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.737917953e-19 lub1 = 1.017341409e-25 wub1 = 1.582997248e-25 pub1 = -3.102278857e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.447139919e-01 lvth0 = -2.195717603e-07 wvth0 = -1.305514161e-07 pvth0 = 2.304181662e-13
+ k1 = 0.64774
+ k2 = 4.910264199e-02 lk2 = -8.312671054e-08 wk2 = -4.507231781e-08 pk2 = 8.723300379e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.889959278e-09 wua = 3.840038595e-18
+ ub = 2.860497637e-18 wub = 1.070410758e-25
+ uc = 4.414740990e-11 wuc = 2.144821557e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.987773017e-03 lu0 = 4.692397691e-10 wu0 = 5.747416245e-10 pu0 = -4.924192753e-16
+ a0 = 2.000068427e+00 la0 = -6.657726332e-07 wa0 = -5.220633599e-07 pa0 = 6.986604698e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 9.917818660e-02 lags = 3.944789433e-07 wags = 1.494571661e-07 pags = -4.139654141e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.854832885e-03 lpdiblc2 = 1.353720531e-08 wpdiblc2 = 1.155768432e-08 ppdiblc2 = -1.420591618e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 6.868625346e-02 ldelta = -3.982300699e-08 wdelta = -4.683489872e-08 pdelta = 4.179018389e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.362938622e+05 lat = -1.885159214e-01 wat = -1.009456466e-01 pat = 1.978282309e-7
+ ute = -1.218144053e-01 wute = -3.404834221e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.592687422e-01 lvth0 = -1.983254636e-07 wvth0 = -2.253401056e-07 pvth0 = 3.687859556e-13
+ k1 = 0.64774
+ k2 = -5.912097746e-02 lk2 = 7.485271795e-08 wk2 = 1.084750902e-08 pk2 = 5.604036574e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.202233871e-09 lua = 4.558428375e-16 wua = 3.315403722e-16 pua = -4.783605620e-22
+ ub = 2.754845221e-18 lub = 1.542261147e-25 wub = 2.179125102e-25 pub = -1.618445763e-31
+ uc = -8.073608746e-11 luc = 1.822986853e-16 wuc = 1.525007079e-16 puc = -1.913038757e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.453452581e-04 lu0 = 3.012748690e-09 wu0 = 2.538745100e-09 pu0 = -3.359373349e-15
+ a0 = 2.021805015e+00 la0 = -6.975026184e-07 wa0 = -5.097641043e-07 pa0 = 6.807066314e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.228024469e-01 lags = 2.140184293e-07 wags = 4.478827735e-08 pags = -2.611750037e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = -1.639628767e+00 lnfactor = 6.097271768e-06 wnfactor = 4.383260695e-06 pnfactor = -6.398464799e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.828704778e-03 lpdiblc2 = 5.240661209e-09 wpdiblc2 = -1.174828784e-08 ppdiblc2 = 1.981497668e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.732044066e-03 ldelta = 5.353415017e-08 wdelta = -2.544854537e-08 pdelta = 1.057145459e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.296557883e-01 lkt1 = -9.005812553e-08 wkt1 = -1.253062194e-08 pkt1 = 1.829157538e-14
+ kt2 = -9.202608700e-02 lkt2 = 5.398314175e-8
+ at = 2.257723765e+05 lat = -2.718218264e-02 wat = 1.674992195e-01 pat = -1.940341623e-7
+ ute = 5.842142473e-01 lute = -1.030625326e-06 wute = -7.657076719e-07 pute = 1.068039706e-12
+ ua1 = 8.009714800e-10 lua1 = -1.531007404e-16
+ ub1 = -3.348293300e-19 lub1 = 3.108527845e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.668850332e-01 lvth0 = 9.342716901e-10 wvth0 = 9.071972059e-08 pvth0 = 6.544753744e-14
+ k1 = 0.64774
+ k2 = 6.768922514e-02 lk2 = -4.685337399e-08 wk2 = -2.993770009e-08 pk2 = 4.474764103e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.375099767e+05 lvsat = -1.319654014e-02 wvsat = 1.529327771e-02 pvsat = -1.467772328e-8
+ ua = -2.704513502e-09 lua = -2.184428689e-17 wua = -1.521695294e-16 pua = -1.411998392e-23
+ ub = 2.954136129e-18 lub = -3.704333489e-26 wub = -6.841668763e-26 pub = 1.129598713e-31
+ uc = 1.462490040e-10 luc = -3.555025625e-17 wuc = -7.821885175e-17 puc = 3.012922168e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.645139086e-03 lu0 = -2.502034365e-10 wu0 = -1.056510003e-09 pu0 = 9.117273614e-17
+ a0 = 8.189900392e-01 la0 = 4.568990548e-07 wa0 = 1.010205856e-06 pa0 = -7.780845376e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 5.508194773e-01 lags = -1.007959156e-07 wags = -3.643776574e-07 pags = 1.315220022e-13
+ b0 = 5.068653630e-07 lb0 = -4.864640321e-13 wb0 = -9.533618939e-13 pb0 = 9.149890777e-19
+ b1 = 2.325991428e-07 lb1 = -2.232370273e-13 wb1 = -7.092873608e-13 pb1 = 6.807385445e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.713350413e+00 wnfactor = -2.283542951e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.938584188e-02 lpdiblc2 = 2.752082236e-08 wpdiblc2 = 8.326858090e-09 ppdiblc2 = 5.478553759e-16
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.288997439e-02 ldelta = 7.314576543e-09 wdelta = -2.098212208e-08 pdelta = 6.284804841e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.818528621e-01 lkt1 = -3.996198396e-08 wkt1 = -1.689367379e-08 pkt1 = 2.247901439e-14
+ kt2 = -2.180719750e-02 lkt2 = -1.340943745e-8
+ at = 3.201167328e+05 lat = -1.177291786e-01 wat = -6.333308374e-02 pat = 2.750714066e-8
+ ute = -4.440801196e-01 lute = -4.371980700e-08 wute = 3.723548224e-07 pute = -2.421577241e-14
+ ua1 = 4.070694500e-10 lua1 = 2.249467329e-16
+ ub1 = 5.630394850e-19 lub1 = -5.508768107e-25 wub1 = -2.869859255e-41 pub1 = 2.736911063e-47
+ uc1 = -2.194613080e-11 luc1 = 1.150272929e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -4.962467785e-01 lvth0 = 6.040833412e-08 wvth0 = 4.285145148e-07 pvth0 = -8.985361922e-14
+ k1 = 0.64774
+ k2 = -1.087877167e-01 lk2 = 3.428190003e-08 wk2 = 9.610472591e-08 pk2 = -1.320036433e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.181905300e+05 lvsat = -4.314424499e-03 wvsat = 9.052395782e-03 pvsat = -1.180847781e-8
+ ua = -2.354576561e-09 lua = -1.827277954e-16 wua = -5.132851588e-16 pua = 1.519029267e-22
+ ub = 2.093061851e-18 lub = 3.588355646e-25 wub = 5.139627657e-25 pub = -1.547890823e-31
+ uc = 1.137836906e-10 luc = -2.062432842e-17 wuc = -5.976079263e-17 puc = 2.164312900e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.535319273e-03 lu0 = -1.997137772e-10 wu0 = -1.714539952e-09 pu0 = 3.937020055e-16
+ a0 = 2.112123481e+00 la0 = -1.376190449e-07 wa0 = -9.963231017e-07 pa0 = 1.444171505e-13
+ keta = -1.176195491e-02 lketa = -3.760962317e-10 wketa = -2.494545072e-09 pketa = 1.146867097e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.315787691e-01 wags = -7.830478701e-8
+ b0 = -1.642697271e-06 lb0 = 5.017973888e-13 wb0 = 3.034996672e-12 pb0 = -9.186587729e-19
+ b1 = -5.551192378e-07 lb1 = 1.389164982e-13 wb1 = 1.692779494e-12 pb1 = -4.236116918e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 4.713350413e+00 wnfactor = -2.283542951e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -8.380581845e-02 lpdiblc2 = 5.713790659e-08 wpdiblc2 = 4.760408645e-08 ppdiblc2 = -1.750985036e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -8.821774543e-03 ldelta = 3.568655312e-08 wdelta = 9.558212866e-08 pdelta = -4.730560944e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.770573649e-01 lkt1 = 3.808286201e-09 wkt1 = 1.746257551e-08 pkt1 = 6.683728776e-15
+ kt2 = -7.233698973e-02 lkt2 = 9.821634527e-09 wkt2 = 9.688746978e-08 pkt2 = -4.454401423e-14
+ at = 1.424300879e+05 lat = -3.603774366e-02 wat = -5.253572802e-03 pat = 8.050855116e-10
+ ute = -6.280372522e-01 lute = 4.085448470e-08 wute = 3.648493470e-07 pute = -2.076513008e-14
+ ua1 = 7.087088751e-10 lua1 = 8.626800716e-17 wua1 = 5.721924709e-16 pua1 = -2.630654885e-22
+ ub1 = -3.120318652e-19 lub1 = -1.485627575e-25 wub1 = -1.211754179e-24 pub1 = 5.571039838e-31
+ uc1 = 3.224846359e-11 luc1 = -1.341323549e-17 wuc1 = -8.896638057e-17 puc1 = 4.090229347e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.868565732e-01 wvth0 = 2.099485795e-8
+ k1 = 0.64774
+ k2 = 1.825397216e-02 wk2 = -2.467105478e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.694093041e-09 wua = -2.017015980e-16
+ ub = 2.757516609e-18 wub = 1.914977057e-25
+ uc = 7.060795191e-11 wuc = -6.319424287e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.964266806e-03 wu0 = -5.640795556e-10
+ a0 = 1.254982334e+00 wa0 = 2.810683114e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.160462985e-01 wags = 2.281646240e-7
+ b0 = -2.317672267e-07 wb0 = 2.432160641e-13
+ b1 = -2.826228170e-07 wb1 = 2.965838189e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.669956697e-03 wpdiblc2 = -1.340875322e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.201855896e-02 wdelta = 9.323282458e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.504878364e-01 wkt1 = -7.436261271e-8
+ kt2 = -0.055045
+ at = 2.636706353e+05 wat = 1.111245810e-2
+ ute = -2.995155341e-01 wute = 8.149135942e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.868565732e-01 wvth0 = 2.099485795e-8
+ k1 = 0.64774
+ k2 = 1.825397216e-02 wk2 = -2.467105478e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.694093041e-09 wua = -2.017015980e-16
+ ub = 2.757516609e-18 wub = 1.914977057e-25
+ uc = 7.060795191e-11 wuc = -6.319424287e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.964266806e-03 wu0 = -5.640795556e-10
+ a0 = 1.254982334e+00 wa0 = 2.810683114e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.160462985e-01 wags = 2.281646240e-7
+ b0 = -2.317672267e-07 wb0 = 2.432160641e-13
+ b1 = -2.826228170e-07 wb1 = 2.965838189e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.669956697e-03 wpdiblc2 = -1.340875322e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.201855896e-02 wdelta = 9.323282458e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.504878364e-01 wkt1 = -7.436261271e-8
+ kt2 = -0.055045
+ at = 2.636706353e+05 wat = 1.111245810e-2
+ ute = -2.995155341e-01 wute = 8.149135942e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.473870848e-01 lvth0 = -3.141672607e-07 wvth0 = -2.656387943e-08 pvth0 = 3.785556599e-13
+ k1 = 0.64774
+ k2 = 5.608266786e-02 lk2 = -3.011069606e-07 wk2 = -3.603219982e-08 pk2 = 2.671697597e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.631805821e-09 lua = -4.957907057e-16 wua = -2.151237613e-16 pua = 1.068370643e-22
+ ub = 2.606521276e-18 lub = 1.201885103e-24 wub = 2.637283164e-25 pub = -5.749376039e-31
+ uc = 6.347964166e-11 luc = 5.673956748e-17 wuc = 1.161010228e-18 puc = -5.954238863e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.826837477e-03 lu0 = 1.093903106e-09 wu0 = -4.360985367e-10 pu0 = -1.018696915e-15
+ a0 = 1.007702303e+00 la0 = 1.968287221e-06 wa0 = 4.497586132e-07 pa0 = -1.342732630e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -2.774021344e-01 lags = 1.284352114e-06 wags = 3.405814684e-07 pags = -8.948099773e-13
+ b0 = -1.632795400e-07 lb0 = -5.451448640e-13 wb0 = 1.713452227e-13 pb0 = 5.720739300e-19
+ b1 = -2.943582889e-07 lb1 = 9.341142260e-14 wb1 = 3.088989997e-13 pb1 = -9.802576005e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.201194122e-03 lpdiblc2 = 3.081339272e-08 wpdiblc2 = -5.894832481e-10 ppdiblc2 = -5.980893059e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -4.572089290e-03 ldelta = 1.320574124e-07 wdelta = 8.219040816e-09 pdelta = -5.800041038e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.802123333e-01 lkt1 = 2.365995638e-07 wkt1 = -7.433493815e-08 pkt1 = -2.202826068e-16
+ kt2 = -0.055045
+ at = 2.517890566e+05 lat = 9.457439664e-02 wat = 2.591834958e-02 pat = -1.178511947e-7
+ ute = -4.152788368e-01 lute = 9.214469487e-07 wute = -3.530546367e-08 pute = 3.458877493e-13
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -2.934552795e-19 lub1 = 1.140833394e-24 wub1 = 6.914628064e-26 pub1 = -5.503871073e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.936522514e-01 lvth0 = -1.309687672e-07 wvth0 = 4.273949232e-08 pvth0 = 1.041316336e-13
+ k1 = 0.64774
+ k2 = -1.750953645e-02 lk2 = -9.700229611e-09 wk2 = 3.282526961e-08 pk2 = -5.488604854e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.884318497e-09 lua = 5.040963646e-16 wua = -1.059632286e-16 pua = -3.254113550e-22
+ ub = 3.074396941e-18 lub = -6.507855606e-25 wub = 8.275024716e-27 pub = 4.365935679e-31
+ uc = 7.780871988e-11 wuc = -1.387589580e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.925877599e-03 lu0 = 7.017289831e-10 wu0 = -6.031143868e-10 pu0 = -3.573559030e-16
+ a0 = 1.750763067e+00 la0 = -9.740476378e-07 wa0 = -3.678089968e-08 pa0 = 5.838422060e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -4.260503108e-02 lags = 3.546142846e-07 wags = 1.207274798e-07 pags = -2.424314594e-14
+ b0 = -3.524277357e-07 lb0 = 2.038347040e-13 wb0 = 3.698369610e-13 pb0 = -2.139037307e-19
+ b1 = -2.619058222e-07 lb1 = -3.509223225e-14 wb1 = 2.748434460e-13 pb1 = 3.682571834e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.447540278e-03 lpdiblc2 = 2.032506669e-08 wpdiblc2 = -1.422332907e-09 ppdiblc2 = -2.683016622e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.405204175e-02 ldelta = -2.088449046e-08 wdelta = -1.340688454e-08 pdelta = 2.763284756e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.204611965e-01 wkt1 = -7.439056858e-8
+ kt2 = -0.055045
+ at = 3.001146598e+05 lat = -9.678291079e-02 wat = 3.319404806e-03 pat = -2.836502311e-8
+ ute = -1.339493575e-01 lute = -1.925474569e-07 wute = 2.289901608e-08 pute = 1.154125606e-13
+ ua1 = 6.9609e-10
+ ub1 = 1.088390903e-19 lub1 = -4.521517372e-25 wub1 = -1.382925613e-25 pub1 = 2.710188470e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.604815752e-01 wvth0 = 9.587465425e-8
+ k1 = 0.64774
+ k2 = -2.245926453e-02 wk2 = 3.002460378e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.627093665e-09 wua = -2.720106097e-16
+ ub = 2.742321135e-18 wub = 2.310552609e-25
+ uc = 7.780871988e-11 wuc = -1.387589580e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.283948263e-03 wu0 = -7.854620857e-10
+ a0 = 1.253736590e+00 wa0 = 2.611357764e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.383437045e-01 wags = 1.083569500e-7
+ b0 = -2.484171711e-07 wb0 = 2.606884825e-13
+ b1 = -2.798123064e-07 wb1 = 2.936344747e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.181879512e-02 wpdiblc2 = -2.791393564e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.339533020e-02 wdelta = 6.933055621e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.204611965e-01 wkt1 = -7.439056858e-8
+ kt2 = -0.055045
+ at = 2.507293245e+05 wat = -1.115439191e-2
+ ute = -2.322003879e-01 wute = 8.179048722e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -6.192292011e-01 lvth0 = 3.777068469e-07 wvth0 = 2.573414800e-07 pvth0 = -2.357011990e-13
+ k1 = 0.64774
+ k2 = -1.237086042e-01 lk2 = 1.477987236e-07 wk2 = 7.862563539e-08 pk2 = -7.094535590e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.632068748e+04 lvsat = 1.130420365e-01 wvsat = 8.126465968e-02 pvsat = -1.186260870e-7
+ ua = -1.827593103e-09 lua = -1.167070946e-15 wua = -1.111004901e-15 pua = 1.224721916e-21
+ ub = 1.881969554e-18 lub = 1.255898219e-24 wub = 1.133906489e-24 pub = -1.317937080e-30
+ uc = 1.248148530e-10 luc = -6.861720286e-17 wuc = -6.320403791e-17 puc = 7.200675545e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 5.276213592e-03 lu0 = -2.908209315e-09 wu0 = -2.740638068e-09 pu0 = 2.854068140e-15
+ a0 = 3.834535850e-01 la0 = 1.270395617e-06 wa0 = 1.209518610e-06 pa0 = -1.384401841e-12
+ keta = -1.064964207e-02 lketa = -2.817839987e-09 wketa = -2.025713750e-09 pketa = 2.957035647e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 5.798021734e-01 lags = -6.444190000e-07 wags = -3.298465217e-07 pags = 6.396675177e-13
+ b0 = 2.265659339e-07 lb0 = -6.933565875e-13 wb0 = -2.377578379e-13 pb0 = 7.276070162e-19
+ b1 = 4.614707060e-07 lb1 = -1.082087877e-12 wb1 = -4.842664360e-13 pb1 = 1.135540854e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 6.589225566e-03 lpdiblc2 = 7.633864163e-09 wpdiblc2 = -1.464517283e-08 ppdiblc2 = 1.730355429e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.080112907e-02 ldelta = 1.229057814e-07 wdelta = 4.332183544e-08 pdelta = -6.222699649e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -2.347183038e-01 lkt1 = -4.171131877e-07 wkt1 = -3.220374283e-07 pkt1 = 3.615025035e-13
+ kt2 = -2.187393836e-01 lkt2 = 2.389528765e-07 wkt2 = 1.329726801e-07 pkt2 = -1.941068697e-13
+ at = 2.789164211e+05 lat = -4.114611415e-02 wat = 1.117299654e-01 pat = -1.793804405e-7
+ ute = -2.225308097e-01 lute = -1.411516677e-08 wute = 8.088897753e-08 pute = 1.315978778e-15
+ ua1 = 1.009910354e-09 lua1 = -4.580992619e-16 wua1 = -2.192600366e-16 pua1 = 3.200648385e-22
+ ub1 = -5.470613180e-19 lub1 = 6.206584290e-25 wub1 = 2.227158238e-25 pub1 = -3.251094238e-31
+ uc1 = 9.220990490e-11 luc1 = -1.491439784e-16 wuc1 = -1.072179433e-16 puc1 = 1.565113927e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -3.576541407e-01 lvth0 = 1.266601828e-07 wvth0 = 8.103284053e-08 pvth0 = -6.648898218e-14
+ k1 = 0.64774
+ k2 = 3.043344871e-02 lk2 = -1.391116839e-10 wk2 = 9.158437180e-09 pk2 = -4.274212413e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.998624180e+05 lvsat = -3.431963944e-02 wvsat = -5.013924951e-02 pvsat = 7.488814879e-9
+ ua = -3.126366219e-09 lua = 7.942655241e-17 wua = 2.905218682e-16 pua = -1.203934001e-22
+ ub = 3.371974735e-18 lub = -1.741342528e-25 wub = -5.068956849e-25 pub = 2.568228064e-31
+ uc = 6.331084342e-11 luc = -9.588729639e-18 wuc = 8.816288089e-18 puc = 2.885247571e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.434693424e-03 lu0 = -1.810603339e-10 wu0 = 2.137292544e-10 pu0 = 1.861410254e-17
+ a0 = 2.207727740e+00 la0 = -4.804515036e-07 wa0 = -4.471327105e-07 pa0 = 2.055692637e-13
+ keta = -1.358565664e-02 wketa = 1.055334071e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.145143683e-01 lags = 2.195130097e-08 wags = 3.338223495e-07 pags = 2.711318581e-15
+ b0 = -1.596017004e-06 lb0 = 1.055867387e-12 wb0 = 1.253398656e-12 pb0 = -7.035304290e-19
+ b1 = -1.842898358e-06 lb1 = 1.129530332e-12 wb1 = 1.468735565e-12 pb1 = -7.388528164e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.609295702e-02 lpdiblc2 = -1.487342103e-09 wpdiblc2 = -2.890452252e-08 ppdiblc2 = 3.098896515e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.875671355e-02 ldelta = 2.735514197e-08 wdelta = -6.150706422e-09 pdelta = -1.474572444e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.659154525e-01 lkt1 = -3.271724239e-09 wkt1 = 7.132144044e-08 pkt1 = -1.602367078e-14
+ kt2 = 6.281688107e-02 lkt2 = -3.127074853e-08 wkt2 = -8.880433880e-08 pkt2 = 1.874362413e-14
+ at = 4.456865844e+05 lat = -2.012037784e-01 wat = -1.951058348e-01 pat = 1.151052187e-7
+ ute = -7.493814870e-02 lute = -1.557672232e-07 wute = -1.502202354e-08 pute = 9.336656205e-14
+ ua1 = -1.397507771e-11 lua1 = 5.245747813e-16 wua1 = 4.418432853e-16 pua1 = -3.144290747e-22
+ ub1 = 1.211546764e-18 lub1 = -1.067165678e-24 wub1 = -6.805422414e-25 pub1 = 5.417925043e-31
+ uc1 = -9.113814615e-11 luc1 = 2.682431357e-17 wuc1 = 7.260996253e-17 puc1 = -1.607843991e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.200118850e-02 lvth0 = -2.765626203e-08 wvth0 = -6.915785883e-08 pvth0 = 2.561191848e-15
+ k1 = 0.64774
+ k2 = -5.242811922e-02 lk2 = 3.795649417e-08 wk2 = 3.696107700e-08 pk2 = -1.705647607e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.904192465e+05 lvsat = -2.997814131e-02 wvsat = -6.674427486e-02 pvsat = 1.512297528e-8
+ ua = -3.090501461e-09 lua = 6.293772985e-17 wua = 2.589929590e-16 pua = -1.058979842e-22
+ ub = 2.660073422e-18 lub = 1.531623757e-25 wub = -8.105804344e-26 pub = 6.104395078e-32
+ uc = 1.431885505e-11 luc = 1.293533702e-17 wuc = 4.461740688e-17 puc = -1.357431679e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.383850168e-03 lu0 = 3.020648534e-10 wu0 = 5.432074239e-10 pu0 = -1.328634859e-16
+ a0 = 1.1627
+ keta = -1.722141262e-02 lketa = 1.671538808e-09 wketa = 3.234598929e-09 pketa = -1.001917018e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -7.847497015e-01 lags = 3.300919954e-07 wags = 1.093168077e-06 pags = -3.463978798e-13
+ b0 = 1.939084068e-06 lb0 = -5.693953306e-13 wb0 = -7.237175015e-13 pb0 = 2.054487245e-19
+ b1 = 9.030021305e-07 lb1 = -1.328974178e-13 wb1 = 1.626298459e-13 pb1 = -1.383707119e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.792390015e-03 lpdiblc2 = 4.167843579e-09 wpdiblc2 = -4.432129831e-08 ppdiblc2 = 3.807682782e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.528726402e-01 ldelta = -2.510965531e-08 wdelta = -7.409966679e-08 pdelta = 1.649381009e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.944366650e-01 lkt1 = 5.581590322e-08 wkt1 = 1.406401783e-07 pkt1 = -4.789296051e-14
+ kt2 = 1.602871186e-01 lkt2 = -7.608269023e-08 wkt2 = -1.472278042e-07 pkt2 = 4.560381236e-14
+ at = -5.965818746e+04 lat = 3.112848044e-02 wat = 2.068174592e-01 pat = -6.967901573e-8
+ ute = -8.296308305e-01 lute = 1.912027372e-07 wute = 5.764012449e-07 pute = -1.785402856e-13
+ ua1 = 1.960985545e-09 lua1 = -3.834133652e-16 wua1 = -7.419441622e-16 pua1 = 2.298172042e-22
+ ub1 = -2.920996469e-18 lub1 = 8.327710739e-25 wub1 = 1.526088059e-24 pub1 = -4.727057762e-31
+ uc1 = -1.624596608e-10 luc1 = 5.961437994e-17 wuc1 = 1.153599358e-16 puc1 = -3.573274011e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -9.079398922e-02 wvth0 = -9.652466279e-8
+ k1 = 0.64774
+ k2 = 5.984653294e-02 wk2 = -2.739760323e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.406118400e-09 wua = 2.250849779e-16
+ ub = 3.775680869e-18 wub = -4.187879157e-25
+ uc = 5.984835477e-11 wuc = 1.298567180e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.614885955e-03 wu0 = 2.447366279e-10
+ a0 = 2.092557968e+00 wa0 = -2.209728485e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.697004740e-01 wags = -2.428104199e-7
+ b0 = 7.434122708e-07 wb0 = -3.413045763e-13
+ b1 = 4.554371000e-08 wb1 = 9.988145895e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 1.516110046e-03 wpdiblc2 = -6.492619474e-10
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.797151477e-03 wdelta = 2.263835451e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.911952308e-01 wkt1 = 1.298567180e-7
+ kt2 = -0.055045
+ at = 2.535045069e+05 wat = 1.720601514e-2
+ ute = -6.782284054e-01 wute = 2.351488736e-7
+ ua1 = 6.8217e-10
+ ub1 = -5.798356185e-20 wub1 = -5.523239074e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 7.436682648e-02 lvth0 = -3.296568591e-06 wvth0 = -1.955217254e-07 pvth0 = 1.975956620e-12
+ k1 = 0.64774
+ k2 = 1.146047477e-01 lk2 = -1.092960276e-06 wk2 = -6.021956762e-08 pk2 = 6.551182037e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.406118400e-09 wua = 2.250849779e-16
+ ub = 3.775680869e-18 wub = -4.187879157e-25
+ uc = 5.984835477e-11 wuc = 1.298567180e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.502653530e-03 lu0 = 2.240131153e-09 wu0 = 3.120085192e-10 pu0 = -1.342730133e-15
+ a0 = 1.688032644e+00 la0 = 8.074224322e-06 wa0 = 2.149882123e-08 pa0 = -4.839673910e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.697004740e-01 wags = -2.428104199e-7
+ b0 = 1.055893114e-06 lb0 = -6.237039509e-12 wb0 = -5.286049687e-13 pb0 = 3.738469008e-18
+ b1 = -1.314989892e-07 lb1 = 3.533728016e-12 wb1 = 2.060004988e-13 pb1 = -2.118109505e-18
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 4.126891095e-03 lpdiblc2 = -5.211053704e-08 wpdiblc2 = -2.214158887e-09 ppdiblc2 = 3.123495168e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.316397107e-02 ldelta = -2.667983774e-07 wdelta = -5.748209480e-09 pdelta = 1.599184138e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.911952308e-01 wkt1 = 1.298567180e-7
+ kt2 = -0.055045
+ at = 2.141776519e+05 lat = 7.849541940e-01 wat = 4.077845337e-02 pat = -4.704999740e-7
+ ute = -6.782284054e-01 wute = 2.351488736e-7
+ ua1 = 6.8217e-10
+ ub1 = 3.138322412e-21 lub1 = -1.219977529e-24 wub1 = -9.186872592e-26 pub1 = 7.312520911e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -5.904819753e-01 lvth0 = 1.995461659e-06 wvth0 = 1.790865117e-07 pvth0 = -1.005831295e-12
+ k1 = 0.64774
+ k2 = -1.182723751e-01 lk2 = 7.606834019e-07 wk2 = 6.847586424e-08 pk2 = -3.692652600e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.472384212e-09 lua = 5.274592941e-16 wua = 2.887172452e-16 pua = -5.064969391e-22
+ ub = 4.176623365e-18 lub = -3.191402030e-24 wub = -6.773877357e-25 pub = 2.058389917e-30
+ uc = 1.060162661e-10 luc = -3.674850325e-16 wuc = -2.433535741e-17 puc = 1.947369881e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.379464306e-03 lu0 = -4.739063428e-09 wu0 = -1.679439531e-10 pu0 = 2.477571559e-15
+ a0 = 3.101515483e+00 la0 = -3.176745702e-06 wa0 = -8.052688190e-07 pa0 = 1.741189814e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.904733903e-01 lags = -9.613222203e-07 wags = -2.995009853e-07 pags = 4.512427275e-13
+ b0 = -2.577757892e-07 lb0 = 4.219436543e-12 wb0 = 2.279860855e-13 pb0 = -2.283806636e-18
+ b1 = 4.960502471e-07 lb1 = -1.461407018e-12 wb1 = -1.648702960e-13 pb1 = 8.339293037e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 2.122913568e-03 lpdiblc2 = -3.615937692e-08 wpdiblc2 = -2.581946749e-09 ppdiblc2 = 3.416245112e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.249104903e-03 ldelta = -3.267764591e-08 wdelta = 9.224240621e-09 pdelta = 4.074145412e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.028106176e+00 lkt1 = 1.089776897e-06 wkt1 = 1.941317354e-07 pkt1 = -5.116130698e-13
+ kt2 = -0.055045
+ at = 3.558881185e+05 lat = -3.430256922e-01 wat = -3.647841994e-02 pat = 1.444454234e-7
+ ute = -1.254849582e+00 lute = 4.589760407e-06 wute = 4.679315616e-07 pute = -1.852892001e-12
+ ua1 = 6.683900700e-10 lua1 = 1.096847978e-16
+ ub1 = -1.780957344e-19 lub1 = 2.226002542e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -7.710606428e-02 lvth0 = -3.737860487e-08 wvth0 = -8.705785916e-08 pvth0 = 4.803387746e-14
+ k1 = 0.64774
+ k2 = 8.473937114e-02 lk2 = -4.319236045e-08 wk2 = -2.846252111e-08 pk2 = 1.458651139e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.293999387e-09 lua = -1.789000171e-16 wua = 1.395986772e-16 pua = 8.397531024e-23
+ ub = 3.280303632e-18 lub = 3.578000342e-25 wub = -1.151450340e-25 pub = -1.679506205e-31
+ uc = 1.321115660e-11 wuc = 2.484375444e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.384669552e-03 lu0 = -7.999248980e-10 wu0 = 3.206826342e-10 pu0 = 5.427324301e-16
+ a0 = 2.060081615e+00 la0 = 9.470720576e-07 wa0 = -2.221858185e-07 pa0 = -5.676730972e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.760153667e-01 lags = 6.798279386e-07 wags = -1.301927493e-07 pags = -2.191755597e-13
+ b0 = 1.163634492e-06 lb0 = -1.408992819e-12 wb0 = -5.388877063e-13 pb0 = 7.528218612e-19
+ b1 = 7.628223154e-08 lb1 = 2.007693815e-13 wb1 = 7.213420299e-14 pb1 = -1.045492612e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -1.923241407e-02 lpdiblc2 = 4.840238170e-08 wpdiblc2 = 1.097319037e-08 ppdiblc2 = -1.951250309e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -5.727314582e-02 ldelta = 1.693648001e-07 wdelta = 4.133325024e-08 pdelta = -8.640219670e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.013426816e-01 lkt1 = -2.041248503e-07 wkt1 = 3.402943181e-08 pkt1 = 1.223520270e-13
+ kt2 = -0.055045
+ at = 3.056525575e+05 lat = -1.441054296e-1
+ ute = -1.499636517e-01 lute = 2.146883463e-07 wute = 3.249795199e-08 pute = -1.286837654e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -9.617921385e-02 wvth0 = -6.254765252e-8
+ k1 = 0.64774
+ k2 = 6.269964135e-02 wk2 = -2.101947409e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.385286549e-09 wua = 1.824486888e-16
+ ub = 3.462877957e-18 wub = -2.008450572e-25
+ uc = 1.321115660e-11 wuc = 2.484375444e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 9.764925405e-04 wu0 = 5.976222592e-10
+ a0 = 2.543343285e+00 wa0 = -5.118518969e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.229106026e-01 wags = -2.420312796e-7
+ b0 = 4.446689000e-07 wb0 = -1.547459223e-13
+ b1 = 1.787286566e-07 wb1 = 1.878593854e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 5.465828918e-03 wpdiblc2 = 1.016561674e-9
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.914848965e-02 wdelta = -2.755126701e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.055012989e-01 wkt1 = 9.646189871e-8
+ kt2 = -0.055045
+ at = 232120.0
+ ute = -4.041480806e-02 wute = -3.316540579e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = 1.140769277e-01 lvth0 = -3.069214026e-07 wvth0 = -1.822007469e-07 pvth0 = 1.746636045e-13
+ k1 = 0.64774
+ k2 = 1.289124583e-01 lk2 = -9.665415953e-08 wk2 = -7.279492425e-08 pk2 = 7.557921337e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.918191587e+05 lvsat = -3.912993570e-01 wvsat = -1.258264330e-01 pvsat = 1.836751356e-7
+ ua = -4.576715022e-09 lua = 1.739187714e-15 wua = 5.368132799e-16 pua = -5.172837118e-22
+ ub = 5.345945005e-18 lub = -2.748807124e-24 wub = -9.423934688e-25 pub = 1.082475294e-30
+ uc = -8.966149132e-11 luc = 1.501683478e-16 wuc = 6.535265394e-17 puc = -5.913286605e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = -2.925385563e-04 lu0 = 1.852468143e-09 wu0 = 5.972608322e-10 pu0 = 5.275930003e-19
+ a0 = 4.686504709e+00 la0 = -3.128479890e-06 wa0 = -1.369721628e-06 pa0 = 1.252275340e-12
+ keta = -7.470874428e-02 lketa = 9.069243446e-08 wketa = 3.637118399e-08 pketa = -5.309283584e-14
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -9.927243005e-01 lags = 2.504398050e-06 wags = 6.127227017e-07 pags = -1.247727124e-12
+ b0 = -8.884610589e-07 lb0 = 1.946036457e-12 wb0 = 4.305871115e-13 pb0 = -8.544398961e-19
+ b1 = -7.779787959e-07 lb1 = 1.396553704e-12 wb1 = 2.586571166e-13 pb1 = -3.501519522e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.291112804e-01 wpclm = 3.351883249e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -4.715720763e-02 lpdiblc2 = 7.681647760e-08 wpdiblc2 = 1.757033173e-08 ppdiblc2 = -2.416436584e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.099183397e-02 ldelta = 1.190667812e-08 wdelta = -5.704703016e-09 pdelta = 4.305644026e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.219923876e+00 lkt1 = 6.049533576e-07 wkt1 = 2.684928215e-07 pkt1 = -2.511221396e-13
+ kt2 = 3.104333000e-03 lkt2 = -8.488348885e-8
+ at = 1.027896501e+06 lat = -1.161634747e+00 wat = -3.372071964e-01 pat = 4.922382050e-7
+ ute = -1.894130284e-01 lute = 2.175001522e-07 wute = 6.103824564e-08 pute = -1.375137802e-13
+ ua1 = 3.433807053e-10 lua1 = 5.148673930e-16 wua1 = 1.802565018e-16 pua1 = -2.631294285e-22
+ ub1 = -4.880210018e-19 lub1 = 5.344743274e-25 wub1 = 1.873271763e-25 pub1 = -2.734508456e-31
+ uc1 = -8.666613950e-11 luc1 = 1.119703274e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -1.591643602e-01 lvth0 = -4.467807657e-08 wvth0 = -3.794153696e-08 pvth0 = 3.621082779e-14
+ k1 = 0.64774
+ k2 = 4.277508293e-02 lk2 = -1.398381352e-08 wk2 = 1.760886314e-09 pk2 = 4.024274178e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.645547492e+05 lvsat = -1.731823399e-01 wvsat = -2.897590342e-02 pvsat = 9.072283980e-8
+ ua = -2.778837784e-09 lua = 1.367503439e-17 wua = 8.221401961e-17 pua = -8.098207174e-23
+ ub = 2.092687198e-18 lub = 3.735070566e-25 wub = 2.599067061e-25 pub = -7.143229913e-32
+ uc = 8.813146605e-11 luc = -2.046844304e-17 wuc = -6.061143475e-18 puc = 9.406526022e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.036812071e-03 lu0 = 5.766238791e-10 wu0 = 1.051616542e-09 pu0 = -4.355402994e-16
+ a0 = 3.418373795e+00 la0 = -1.911391245e-06 wa0 = -1.172791534e-06 pa0 = 1.063271682e-12
+ keta = 4.634785522e-02 lketa = -2.549163690e-08 wketa = -3.486869307e-08 pketa = 1.527963618e-14
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.489515562e+00 lags = 1.220683421e-07 wags = -6.276299824e-07 pags = -5.729863566e-14
+ b0 = 1.664343631e-06 lb0 = -5.040178438e-13 wb0 = -7.008549878e-13 pb0 = 2.314616587e-19
+ b1 = 3.726066137e-07 lb1 = 2.922793569e-13 wb1 = 1.407663164e-13 pb1 = -2.370062567e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -9.344276432e-01 lpclm = 3.890023792e-07 wpclm = 5.781341421e-07 ppclm = -2.331672481e-13
+ pdiblc1 = 0.0
+ pdiblc2 = -1.273572964e-01 lpdiblc2 = 1.537885128e-07 wpdiblc2 = 5.707927250e-08 ppdiblc2 = -6.208307174e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.972205229e-02 ldelta = -6.365464891e-08 wdelta = -4.269320853e-08 pdelta = 3.980536220e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -4.563438738e-01 lkt1 = -1.278925500e-07 wkt1 = -5.429534466e-08 pkt1 = 5.867380292e-14
+ kt2 = -0.085339
+ at = -3.552405265e+05 lat = 1.658310149e-01 wat = 2.849682736e-01 pat = -1.048947024e-7
+ ute = 1.633719963e-01 lute = -1.210852753e-07 wute = -1.578646478e-07 pute = 7.257827184e-14
+ ua1 = 9.278490842e-10 lua1 = -4.607613370e-17 wua1 = -1.226842337e-16 pua1 = 2.761794239e-23
+ ub1 = 9.513846034e-19 lub1 = -8.469952022e-25 wub1 = -5.246015628e-25 pub1 = 4.098227617e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.0125e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -2.4699e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = -2.690632801e-02 lvth0 = -1.054837069e-07 wvth0 = -6.621772801e-08 pvth0 = 4.921080662e-14
+ k1 = 0.64774
+ k2 = 6.313987534e-02 lk2 = -2.334652683e-08 wk2 = -3.231014780e-08 pk2 = 1.968843211e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -6.617423650e+05 lvsat = 2.067077584e-01 wvsat = 4.440396907e-01 pvsat = -1.267460796e-7
+ ua = -2.061790088e-09 lua = -3.159876438e-16 wua = -3.576145801e-16 pua = 1.212291270e-22
+ ub = 1.317011342e-18 lub = 7.301240316e-25 wub = 7.239706815e-25 pub = -2.847857118e-31
+ uc = 7.453845146e-11 luc = -1.421905458e-17 wuc = 8.521901228e-18 puc = 2.701971220e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.699113389e-03 lu0 = 2.721308479e-10 wu0 = 3.542392793e-10 pu0 = -1.149211029e-16
+ a0 = -7.390840508e-01 wa0 = 1.139925556e-6
+ keta = -9.098880846e-03 wketa = -1.634030369e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.240346405e+00 lags = -1.142626138e-06 wags = -1.918864479e-06 pags = 5.363464239e-13
+ b0 = 1.741094271e-06 lb0 = -5.393039504e-13 wb0 = -6.050428131e-13 pb0 = 1.874120114e-19
+ b1 = 3.090568317e-06 lb1 = -9.573035363e-13 wb1 = -1.148592951e-12 pb1 = 3.557766667e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = -0.1819
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = 2.5373
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.831045088e-02 wpclm = 7.097318924e-8
+ pdiblc1 = 0.0
+ pdiblc2 = -4.564133840e-02 lpdiblc2 = 1.162196011e-07 wpdiblc2 = -1.469082037e-08 ppdiblc2 = -2.908677155e-14
+ pdiblcb = -0.025
+ drout = 4.663735585e-01 wdrout = -1.882922411e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.249506561e-01 ldelta = -7.525349952e-08 wdelta = -5.736328537e-08 pdelta = 4.654993002e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.347495730e-01 lkt1 = 9.205447025e-08 wkt1 = 2.247434548e-07 pkt1 = -6.961428511e-14
+ kt2 = -0.085339
+ at = -5.123944135e+03 lat = 4.864916196e-03 wat = 1.741297428e-01 pat = -5.393668784e-8
+ ute = 1.320027500e-01 lute = -1.066632643e-07 pute = 2.524354897e-29
+ ua1 = 1.043337168e-09 lua1 = -9.917178040e-17 wua1 = -1.919075604e-16 pua1 = 5.944336683e-23
+ ub1 = -2.250590322e-18 lub1 = 6.251127698e-25 wub1 = 1.124247955e-24 pub1 = -3.482358040e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 1.0e-11
+ cgso = 1.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 3.417e-8
+ dwc = -3.2175e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006926438503
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.29052224e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.164485778e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = 0
+ kvth0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 0
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.109639
+ k1 = 0.43657182
+ k2 = 0.027786788
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.22271988
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.2497576
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.019607598
+ ua = -2.7648397e-10
+ ub = 2.34385173e-18
+ uc = -7.7670696e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200000.0
+ a0 = 1.5017417
+ ags = 0.38244371
+ a1 = 0.0
+ a2 = 1.0
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.013169082
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.075489662
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 746475130.0
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1154444600.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.44169
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.109639
+ k1 = 0.43657182
+ k2 = 0.027786788
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.22271988
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.2497576
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.019607598
+ ua = -2.7648397e-10
+ ub = 2.34385173e-18
+ uc = -7.7670696e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200000.0
+ a0 = 1.5017417
+ ags = 0.38244371
+ a1 = 0.0
+ a2 = 1.0
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.013169082
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.075489662
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 746475130.0
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1154444600.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.44169
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108748660e+00 lvth0 = -7.112810250e-09 wvth0 = -8.907461576e-08 pvth0 = 7.116055256e-13
+ k1 = 4.360518078e-01 lk1 = 4.154309705e-09 wk1 = 5.202494200e-08 pk1 = -4.156204984e-13
+ k2 = 2.819103967e-02 lk2 = -3.229514006e-09 wk2 = -4.044360936e-08 pk2 = 3.230987375e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.235312098e-01 lvoff = 6.481607941e-09 wvoff = 8.116999000e-08 pvoff = -6.484564980e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.201405605e+00 lnfactor = 3.862778035e-07 wnfactor = 4.837405429e-06 pnfactor = -3.864540311e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.932502699e-02 lu0 = 2.257423098e-09 wu0 = 2.826999288e-08 pu0 = -2.258452980e-13
+ ua = -3.021630050e-10 lua = 2.051464722e-16 wua = 2.569075027e-15 pua = -2.052400641e-20
+ ub = 2.324401486e-18 lub = 1.553854689e-25 wub = 1.945911736e-24 pub = -1.554563589e-29
+ uc = -7.712273168e-11 luc = -4.377615734e-18 wuc = -5.482143144e-17 puc = 4.379612890e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.943880576e+05 lvsat = 4.483307809e-02 wvsat = 5.614502657e-01 pvsat = -4.485353184e-6
+ a0 = 1.524697852e+00 la0 = -1.833937180e-07 wa0 = -2.296662555e-06 pa0 = 1.834773858e-11
+ ags = 4.014098279e-01 lags = -1.515178505e-07 wags = -1.897477064e-06 pags = 1.515869759e-11
+ a1 = 0.0
+ a2 = 9.848810403e-01 la2 = 1.207035148e-07 wa2 = 1.511585270e-06 pa2 = -1.207585822e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.635811733e-02 lketa = 2.547678869e-08 wketa = 3.190490233e-07 pketa = -2.548841171e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.175946087e-01 lpclm = -3.363709457e-07 wpclm = -4.212415583e-06 ppclm = 3.365244048e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.389656634e-03 lpdiblc2 = 1.900893826e-09 wpdiblc2 = 2.380513203e-08 ppdiblc2 = -1.901761051e-13
+ pdiblcb = -1.467644794e-04 lpdiblcb = 4.075956659e-10 wpdiblcb = 5.104371697e-09 ppdiblcb = -4.077816192e-14
+ drout = 0.56
+ pscbe1 = 7.505188577e+08 lpscbe1 = -3.230481493e+01 wpscbe1 = -4.045572532e+02 ppscbe1 = 3.231955303e-3
+ pscbe2 = 9.463108264e-09 lpscbe2 = 3.346077183e-16 wpscbe2 = 4.190334466e-15 ppscbe2 = -3.347603731e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.831979289e+00 lbeta0 = -3.162808702e-07 wbeta0 = -3.960825046e-06 pbeta0 = 3.164251638e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.034252636e-10 lagidl = -2.736398594e-17 wagidl = -3.426826314e-16 pagidl = 2.737646994e-21
+ bgidl = 1.142776530e+09 lbgidl = 9.321469104e+01 wbgidl = 1.167339279e+03 pbgidl = -9.325721745e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.425036582e-01 lkt1 = 6.500209282e-09 wkt1 = 8.140293693e-08 pkt1 = -6.503174808e-13
+ kt2 = -3.814118335e-02 lkt2 = 1.439461387e-09 wkt2 = 1.802655567e-08 pkt2 = -1.440118098e-13
+ at = 1.983225665e+04 lat = -1.584373202e-01 wat = -1.984130453e+00 pat = 1.585096025e-5
+ ute = -3.004779279e-01 lute = -1.454550081e-09 wute = -1.821551328e-08 pute = 1.455213676e-13
+ ua1 = 2.227223445e-09 lua1 = -1.248136750e-16 wua1 = -1.563057322e-15 pua1 = 1.248706175e-20
+ ub1 = -8.067528284e-19 lub1 = 1.051561247e-25 wub1 = 1.316883352e-24 pub1 = -1.052040991e-29
+ uc1 = 1.211396142e-10 luc1 = -1.030256012e-17 wuc1 = -1.290202538e-16 puc1 = 1.030726035e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.122759258e+00 lvth0 = 4.877364531e-08 wvth0 = 1.401481030e-07 pvth0 = -2.027341004e-13
+ k1 = 4.493657172e-01 lk1 = -4.895314383e-08 wk1 = -5.951765964e-07 pk1 = 2.165982302e-12
+ k2 = 1.965123111e-02 lk2 = 3.083467214e-08 wk2 = 2.815734565e-07 pk2 = -9.613854759e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.442199869e-01 ldsub = 6.294442095e-08 wdsub = 1.578721228e-06 pdsub = -6.297313746e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.097347255e-01 lvoff = -4.855077438e-08 wvoff = -2.306790003e-07 pvoff = 5.954685840e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.002861472e+00 lnfactor = -2.810625461e-06 wnfactor = -1.167067584e-05 pnfactor = 2.720318701e-11
+ eta0 = 7.401064685e-02 leta0 = 2.389075108e-08 weta0 = 5.992085608e-07 peta0 = -2.390165052e-12
+ etab = -6.476402461e-02 letab = -2.088562516e-08 wetab = -5.238364148e-07 petab = 2.089515360e-12
+ u0 = 2.366069310e-02 lu0 = -1.503698541e-08 wu0 = -3.338058468e-08 pu0 = 2.007084129e-14
+ ua = 9.272450516e-11 lua = -1.370008470e-15 wua = -3.121327775e-15 pua = 2.174270613e-21
+ ub = 2.623200850e-18 lub = -1.036486351e-24 wub = -2.333901187e-24 pub = 1.525981486e-30
+ uc = -8.615807197e-11 luc = 3.166318211e-17 wuc = 1.275182190e-16 puc = -2.893678725e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.799149686e+05 lvsat = -2.963226514e-01 wvsat = -6.048539334e-01 pvsat = 1.668826468e-7
+ a0 = 1.149595481e+00 la0 = 1.312840879e-06 wa0 = 5.000049791e-06 pa0 = -1.075789839e-11
+ ags = 1.073348097e-01 lags = 1.021509168e-06 wags = 2.547224328e-06 pags = -2.570638448e-12
+ a1 = 0.0
+ a2 = 1.229084975e+00 la2 = -8.533942343e-07 wa2 = -3.023170540e-06 pa2 = 6.012693192e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.501192289e-02 lketa = -1.794316236e-07 wketa = -6.207023588e-07 pketa = 1.199704925e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.647293317e-01 lpclm = 2.385330551e-06 wpclm = 8.603689119e-06 ppclm = -1.746933508e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 7.217847004e-03 lpdiblc2 = -1.336925990e-08 wpdiblc2 = -4.584503763e-08 ppdiblc2 = 8.764936711e-14
+ pdiblcb = 6.199588191e-04 lpdiblcb = -2.650763898e-09 wpdiblcb = -4.414829700e-09 ppdiblcb = -2.807305045e-15
+ drout = 0.56
+ pscbe1 = 6.851606705e+08 lpscbe1 = 2.284004973e+02 wpscbe1 = 8.091145064e+02 ppscbe1 = -1.609223568e-3
+ pscbe2 = 1.011912642e-08 lpscbe2 = -2.282163411e-15 wpscbe2 = -6.284641909e-15 ppscbe2 = 8.307281707e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.340918808e+00 lbeta0 = 1.642495549e-06 wbeta0 = -6.968142227e-06 pbeta0 = 4.363831367e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.504514984e-11 lagidl = 2.055066986e-16 wagidl = 9.873101499e-16 pagidl = -2.567521312e-21
+ bgidl = 1.331365855e+09 lbgidl = -6.590436080e+02 wbgidl = -2.334678558e+03 pbgidl = 4.643372143e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.277110086e-01 lkt1 = -5.250574678e-08 wkt1 = -3.270417800e-07 pkt1 = 9.789153974e-13
+ kt2 = -3.548113669e-02 lkt2 = -9.171118947e-09 wkt2 = -1.081851686e-08 pkt2 = -2.895256535e-14
+ at = -3.136423608e+05 lat = 1.171749577e+00 wat = 5.261722303e+00 pat = -1.305180443e-5
+ ute = -2.935034937e-01 lute = -2.927466138e-08 wute = -9.557452919e-07 pute = 3.885205776e-12
+ ua1 = 1.930766960e-09 lua1 = 1.057712705e-15 wua1 = 7.521818200e-15 pua1 = -2.375132567e-20
+ ub1 = -5.690430214e-19 lub1 = -8.430373928e-25 wub1 = -5.130996646e-24 pub1 = 1.519934518e-29
+ uc1 = 8.453246673e-11 luc1 = 1.357185922e-16 wuc1 = 1.835089605e-15 puc1 = -6.803852856e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.096635140e+00 lvth0 = -3.183830430e-09 wvth0 = -1.219416244e-07 pvth0 = 3.185282958e-13
+ k1 = 4.209874975e-01 lk1 = 7.487445918e-09 wk1 = 8.705142160e-07 pk1 = -7.490861840e-13
+ k2 = 3.664638724e-02 lk2 = -2.966484037e-09 wk2 = -3.510315989e-07 pk2 = 2.967837406e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.245231430e-01 ldsub = -9.676811721e-08 wdsub = -6.455257977e-06 pdsub = 9.681226476e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.343090447e-01 lvoff = 3.243519242e-10 wvoff = 8.503724761e-08 pvoff = -3.244999001e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.571212030e+00 lnfactor = 3.673916402e-08 wnfactor = 3.855114951e-06 pnfactor = -3.675592516e-12
+ eta0 = 1.024505933e-01 leta0 = -3.267260519e-08 weta0 = -2.246083570e-06 peta0 = 3.268751109e-12
+ etab = -7.530273474e-02 letab = 7.449926597e-11 wetab = 5.305153957e-07 petab = -7.453325403e-15
+ u0 = 1.600368364e-02 lu0 = 1.918110102e-10 wu0 = -1.364038390e-08 pu0 = -1.918985182e-14
+ ua = -5.894234371e-10 lua = -1.330489245e-17 wua = -2.697381327e-15 pua = 1.331096241e-21
+ ub = 2.074848117e-18 lub = 5.411594944e-26 wub = 1.155540208e-24 pub = -5.414063822e-30
+ uc = -6.957681104e-11 luc = -1.314790313e-18 wuc = -8.411295202e-17 puc = 1.315390146e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.333042000e+05 lvsat = -4.732892029e-03 wvsat = -7.590231250e-01 pvsat = 4.735051269e-7
+ a0 = 1.811685334e+00 la0 = -3.969767887e-09 wa0 = -6.086909959e-07 pa0 = 3.971578974e-13
+ ags = 6.300862175e-01 lags = -1.817542500e-08 wags = 3.404384909e-07 pags = 1.818371699e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.402520275e-02 lketa = -2.348355581e-09 wketa = -1.356217703e-07 pketa = 2.349426948e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.430702329e-01 lpclm = -1.682576948e-08 wpclm = -1.026241271e-06 ppclm = 1.683344573e-12
+ pdiblc1 = 3.865953011e-01 lpdiblc1 = 6.771503502e-09 wpdiblc1 = 3.406252192e-07 ppdiblc1 = -6.774592797e-13
+ pdiblc2 = 5.097534716e-04 lpdiblc2 = -2.773391177e-11 wpdiblc2 = -3.170196810e-09 ppdiblc2 = 2.774656454e-15
+ pdiblcb = -6.978912554e-04 lpdiblcb = -2.973142036e-11 wpdiblcb = -7.321909342e-09 ppdiblcb = 2.974498443e-15
+ drout = 5.816813724e-01 ldrout = -4.312143120e-08 wdrout = -2.169126392e-06 pdrout = 4.314110406e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 9.004001941e-09 lpscbe2 = -6.432579521e-17 wpscbe2 = -5.343520813e-15 ppscbe2 = 6.435514193e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.280633849e+00 lbeta0 = -2.264755038e-07 wbeta0 = 3.580778026e-06 pbeta0 = 2.265788264e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.479781125e-10 lagidl = 7.864172316e-19 wagidl = -2.640756676e-16 pagidl = -7.867760109e-23
+ bgidl = 1.009479675e+09 lbgidl = -1.885384214e+01 wbgidl = -9.484000280e+02 pbgidl = 1.886244364e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.571230211e-01 lkt1 = 5.990922543e-09 wkt1 = 4.665148474e-07 pkt1 = -5.993655721e-13
+ kt2 = -4.035397695e-02 lkt2 = 5.203268623e-10 wkt2 = 7.980590052e-10 pkt2 = -5.205642458e-14
+ at = 2.796698942e+05 lat = -8.271367424e-03 wat = -1.716772285e+00 pat = 8.275140987e-7
+ ute = -4.014196268e-01 lute = 1.853564981e-07 wute = 1.032166948e-05 pute = -1.854410615e-11
+ ua1 = 2.276780712e-09 lua1 = 3.695363340e-16 wua1 = 1.416838973e-14 pua1 = -3.697049238e-20
+ ub1 = -8.879763809e-19 lub1 = -2.087204022e-25 wub1 = -7.988004532e-24 pub1 = 2.088156246e-29
+ uc1 = 1.581711189e-10 luc1 = -1.073911389e-17 wuc1 = -2.126081405e-15 puc1 = 1.074401329e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.103462676e+00 lvth0 = 3.567715066e-09 wvth0 = 6.794160859e-08 pvth0 = 1.307584631e-13
+ k1 = 3.626009089e-01 lk1 = 6.522419181e-08 wk1 = 3.379529178e-07 pk1 = -2.224522931e-13
+ k2 = 6.088486525e-02 lk2 = -2.693518778e-08 wk2 = -1.714622965e-07 pk2 = 1.192130445e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.469753064e-01 ldsub = -2.178573881e-07 wdsub = 1.782716347e-06 pdsub = 1.534940806e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.434787499e-01 lvoff = 9.391998282e-09 wvoff = 1.155165391e-07 pvoff = -6.259004695e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.392932729e+00 lnfactor = 2.130342168e-07 wnfactor = -4.211325382e-06 pnfactor = 4.301068337e-12
+ eta0 = 1.378002277e-01 leta0 = -6.762879820e-08 weta0 = 1.993919478e-06 peta0 = -9.240607050e-13
+ etab = -1.483283986e-01 letab = 7.228738745e-08 wetab = 1.038020206e-06 petab = -5.093096073e-13
+ u0 = 1.923299871e-02 lu0 = -3.001561782e-09 wu0 = -3.615455914e-08 pu0 = 3.073740640e-15
+ ua = -3.329492658e-10 lua = -2.669245063e-16 wua = -2.182009776e-15 pua = 8.214607756e-22
+ ub = 2.323395052e-18 lub = -1.916646575e-25 wub = -3.491645699e-24 pub = -8.186010938e-31
+ uc = -6.477667493e-11 luc = -6.061500909e-18 wuc = -3.323576763e-16 puc = 3.770207751e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.974570296e+05 lvsat = -6.817170060e-02 wvsat = -4.539804450e-01 pvsat = 1.718575719e-7
+ a0 = 1.812994089e+00 la0 = -5.263955862e-09 wa0 = 4.538881060e-06 pa0 = -4.693121682e-12
+ ags = 4.386333933e-01 lags = 1.711465293e-07 wags = 3.301312849e-06 pags = -1.109548128e-12
+ a1 = 0.0
+ a2 = 8.148138538e-01 la2 = -1.464897560e-08 wa2 = -1.482061217e-06 pa2 = 1.465565876e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.314527244e-02 lketa = -3.218492269e-09 wketa = 2.107756890e-09 pketa = 9.874609720e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.633949386e-01 lpclm = -3.692426118e-08 wpclm = -7.384055170e-07 ppclm = 1.398712431e-12
+ pdiblc1 = 3.720535046e-01 lpdiblc1 = 2.115144982e-08 wpdiblc1 = 1.795468297e-06 ppdiblc1 = -2.116109954e-12
+ pdiblc2 = 7.537206750e-04 lpdiblc2 = -2.689857602e-10 wpdiblc2 = -4.668789910e-09 ppdiblc2 = 4.256570213e-15
+ pdiblcb = -1.671969296e-03 lpdiblcb = 9.335051313e-10 wpdiblcb = 1.653242344e-07 ppdiblcb = -1.677500937e-13
+ drout = 5.457651998e-01 ldrout = -7.605005539e-09 wdrout = 1.424129443e-06 pdrout = 7.608475095e-13
+ pscbe1 = 7.969604563e+08 lpscbe1 = 3.005713570e+00 wpscbe1 = 3.040930392e+02 ppscbe1 = -3.007084837e-4
+ pscbe2 = 9.233762175e-09 lpscbe2 = -2.915287980e-16 wpscbe2 = -1.127610960e-15 ppscbe2 = 2.266527416e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.992863204e+00 lbeta0 = 2.035832253e-06 wbeta0 = 3.922123529e-05 pbeta0 = -1.258589633e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.909095767e-10 lagidl = -4.166721980e-17 wagidl = -6.405145136e-16 pagidl = 2.935714805e-22
+ bgidl = 9.935672924e+08 lbgidl = -3.118563934e+00 wbgidl = 6.435642293e+02 pbgidl = 3.119986685e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.754280130e-01 lkt1 = 2.409217992e-08 wkt1 = 1.663817167e-07 pkt1 = -3.025729233e-13
+ kt2 = -3.523070398e-02 lkt2 = -4.545924082e-09 wkt2 = -1.842662778e-07 pkt2 = 1.309481461e-13
+ at = 4.439247213e+05 lat = -1.706980384e-01 wat = -1.363097581e+00 pat = 4.777757946e-7
+ ute = -2.560929686e-01 lute = 4.164732565e-08 wute = -1.709417433e-05 pute = 8.566599321e-12
+ ua1 = 3.501774071e-09 lua1 = -8.418228484e-16 wua1 = -5.133902149e-14 pua1 = 2.780782134e-20
+ ub1 = -1.658531144e-18 lub1 = 5.532580868e-25 wub1 = 3.669336537e-23 pub1 = -2.330250380e-29
+ uc1 = 3.529363748e-10 luc1 = -2.033366325e-16 wuc1 = -1.144416457e-15 puc1 = 1.036623125e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.096961525e+00 lvth0 = 3.894973997e-10 wvth0 = 4.151217848e-07 pvth0 = -3.896750962e-14
+ k1 = 5.154033531e-01 lk1 = -9.476339101e-09 wk1 = -2.056382044e-06 pk1 = 9.480662397e-13
+ k2 = -7.801580673e-04 lk2 = 3.210992167e-09 wk2 = 7.295108724e-07 pk2 = -3.212457086e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.784316906e-01 ldsub = 1.119952944e-08 wdsub = 7.214435814e-06 pdsub = -1.120463889e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.267427690e-01 lvoff = 1.210279319e-09 wvoff = 2.351661397e-07 pvoff = -1.210831472e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.805106377e+00 lnfactor = 1.153488555e-08 wnfactor = 6.947230341e-06 pnfactor = -1.154014800e-12
+ eta0 = 3.390588200e-02 leta0 = -1.683796940e-08 weta0 = -3.342112243e-06 peta0 = 1.684565122e-12
+ etab = -4.349753485e-04 letab = -1.327035823e-11 wetab = -6.505431706e-09 petab = 1.327641243e-15
+ u0 = 1.283779815e-02 lu0 = 1.248599159e-10 wu0 = -4.314952314e-09 pu0 = -1.249168795e-14
+ ua = -9.427720475e-10 lua = 3.119955704e-17 wua = 5.883201561e-15 pua = -3.121379091e-21
+ ub = 1.974182722e-18 lub = -2.094522568e-26 wub = -9.452492600e-24 pub = 2.095478131e-30
+ uc = -7.609646532e-11 luc = -5.275949820e-19 wuc = 3.308804176e-16 puc = 5.278356814e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.992219728e+04 lvsat = -9.350471346e-04 wvsat = -2.937943020e-01 pvsat = 9.354737218e-8
+ a0 = 1.780369366e+00 la0 = 1.068529245e-08 wa0 = -2.874347309e-06 pa0 = -1.069016729e-12
+ ags = 8.879649710e-01 lags = -4.851819906e-08 wags = -8.897393415e-06 pags = 4.854033404e-12
+ a1 = 0.0
+ a2 = 7.703722924e-01 la2 = 7.077170512e-09 wa2 = 2.964122434e-06 pa2 = -7.080399259e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.383587559e-02 lketa = 2.007822894e-09 wketa = 6.149905017e-07 pketa = -2.008738903e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.757783535e-01 lpclm = 5.908858790e-09 wpclm = 3.331936055e-06 ppclm = -5.911554530e-13
+ pdiblc1 = 4.384124393e-01 lpdiblc1 = -1.128944260e-08 wpdiblc1 = -4.843452603e-06 ppdiblc1 = 1.129459307e-12
+ pdiblc2 = 7.604466525e-04 lpdiblc2 = -2.722738888e-10 wpdiblc2 = -5.168177975e-08 ppdiblc2 = 2.723981056e-14
+ pdiblcb = 2.375467952e-04 wpdiblcb = -1.778142149e-7
+ drout = 5.018998453e-01 ldrout = 1.383945029e-08 wdrout = 5.812666112e-06 pdrout = -1.384576412e-12
+ pscbe1 = 8.060790874e+08 lpscbe1 = -1.452111603e+00 wpscbe1 = -6.081860784e+02 ppscbe1 = 1.452774086e-4
+ pscbe2 = 8.048535097e-09 lpscbe2 = 2.878931638e-16 wpscbe2 = 6.242502687e-14 ppscbe2 = -2.880245064e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.235084956e-09 lalpha0 = -5.549089824e-16 walpha0 = -1.135602804e-13 palpha0 = 5.551621430e-20
+ alpha1 = 9.276134311e-11 lalpha1 = 3.538762194e-18 walpha1 = 7.241959311e-16 palpha1 = -3.540376648e-22
+ beta0 = 7.705846421e+00 lbeta0 = -2.682038519e-07 wbeta0 = -4.141066586e-05 pbeta0 = 2.683262118e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056778795e-10 wagidl = -4.000419274e-17
+ bgidl = 9.924854795e+08 lbgidl = -2.589698023e+00 wbgidl = 7.517948818e+02 pbgidl = 2.590879495e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.266178953e-01 lkt1 = 2.303776654e-10 wkt1 = -4.053953333e-07 pkt1 = -2.304827683e-14
+ kt2 = -4.494262190e-02 lkt2 = 2.019412340e-10 wkt2 = 1.249191549e-07 pkt2 = -2.020333636e-14
+ at = 9.513885628e+04 lat = -1.870925171e-04 wat = -4.240790133e-01 pat = 1.871778724e-8
+ ute = -1.665587714e-01 lute = -2.123257317e-09 wute = -5.425330174e-09 pute = 2.124225989e-13
+ ua1 = 1.681101245e-09 lua1 = 4.824947608e-17 wua1 = 1.541690583e-14 pua1 = -4.827148846e-21
+ ub1 = -4.297318726e-19 lub1 = -4.746501319e-26 wub1 = -2.068624591e-23 pub1 = 4.748666767e-30
+ uc1 = -5.422306194e-11 luc1 = -4.288598690e-18 wuc1 = -1.810019196e-15 puc1 = 4.290555235e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.111694797e+00 lvth0 = 3.908834132e-09 wvth0 = 1.889121167e-06 pvth0 = -3.910617421e-13
+ k1 = 5.190311829e-01 lk1 = -1.034291882e-08 wk1 = -2.419330537e-06 pk1 = 1.034763746e-12
+ k2 = -2.503657329e-03 lk2 = 3.622684435e-09 wk2 = 9.019394281e-07 pk2 = -3.624337176e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.036552333e-01 ldsub = 5.174381798e-09 wdsub = 4.690930795e-06 pdsub = -5.176742454e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.280998913e-01 lvoff = 1.534455130e-09 wvoff = 3.709402877e-07 pvoff = -1.535155179e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.847221791e+00 lnfactor = 1.474776644e-09 wnfactor = 2.733767566e-06 pnfactor = -1.475449466e-13
+ eta0 = -3.658421472e-02 weta0 = 3.710113328e-6
+ etab = -4.905300834e-04 letab = 1.309705708e-18 wetab = -9.474236925e-10 petab = -1.310303216e-22
+ u0 = 1.302528849e-02 lu0 = 8.007409696e-11 wu0 = -2.307254059e-08 pu0 = -8.011062836e-15
+ ua = -8.720118943e-10 lua = 1.429707924e-17 wua = -1.196041982e-15 pua = -1.430360186e-21
+ ub = 1.900026297e-18 lub = -3.231480537e-27 wub = -2.033466978e-24 pub = 3.232954803e-31
+ uc = -8.030829580e-11 luc = 4.784849643e-19 wuc = 7.522556176e-16 puc = -4.787032587e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.622431241e+04 lvsat = -5.173337526e-05 wvsat = 7.616289011e-02 pvsat = 5.175697706e-9
+ a0 = 1.792752791e+00 la0 = 7.727263646e-09 wa0 = -4.113254795e-06 pa0 = -7.730788978e-13
+ ags = 4.918140472e-01 lags = 4.611037211e-08 wags = 3.073577216e-05 pags = -4.613140858e-12
+ a1 = 0.0
+ a2 = 7.862174314e-01 la2 = 3.292242150e-09 wa2 = 1.378885644e-06 pa2 = -3.293744137e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.556141279e-02 lketa = 3.130196629e-11 wketa = -2.128332752e-07 pketa = -3.131624688e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.970489189e-01 lpclm = 8.279588369e-10 wpclm = 1.203909110e-06 ppclm = -8.283365683e-14
+ pdiblc1 = 3.971394206e-01 lpdiblc1 = -1.430556614e-09 wpdiblc1 = -7.142677733e-07 ppdiblc1 = 1.431209262e-13
+ pdiblc2 = -2.576915399e-04 lpdiblc2 = -2.907121879e-11 wpdiblc2 = 5.017848898e-08 ppdiblc2 = 2.908448166e-15
+ pdiblcb = -2.724839315e-02 lpdiblcb = 6.565566475e-09 wpdiblcb = 2.572033743e-06 ppdiblcb = -6.568561818e-13
+ drout = 5.640284291e-01 ldrout = -1.001204524e-09 wdrout = -4.030266976e-07 pdrout = 1.001661294e-13
+ pscbe1 = 7.999813105e+08 lpscbe1 = 4.464350172e-03 wpscbe1 = 1.869798174e+00 ppscbe1 = -4.466386898e-7
+ pscbe2 = 1.076745325e-08 lpscbe2 = -3.615748147e-16 wpscbe2 = -2.095908306e-13 ppscbe2 = 3.617397723e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.319903354e-09 lalpha0 = 5.540107511e-17 walpha0 = 1.420551142e-13 palpha0 = -5.542635018e-21
+ alpha1 = 1.075759376e-10 walpha1 = -7.579393929e-16
+ beta0 = 6.498208410e+00 lbeta0 = 2.026463977e-08 wbeta0 = 7.940823008e-05 pbeta0 = -2.027388490e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056778795e-10 wagidl = -4.000419274e-17
+ bgidl = 1.009965861e+09 lbgidl = -6.765236785e+00 wbgidl = -9.970407720e+02 pbgidl = 6.768323221e-4
+ cgidl = 2.541335236e+02 lcgidl = 1.095612521e-05 wcgidl = 4.588740156e-03 pcgidl = -1.096112361e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.294555033e-01 lkt1 = 9.081970836e-10 wkt1 = -1.215050779e-07 pkt1 = -9.086114213e-14
+ kt2 = -4.678647856e-02 lkt2 = 6.423832743e-10 wkt2 = 3.093889413e-07 pkt2 = -6.426763424e-14
+ at = 9.211512097e+04 lat = 5.351871368e-04 wat = -1.215675333e-01 pat = -5.354312999e-8
+ ute = -1.968199601e-01 lute = 5.105232829e-09 wute = 3.022074116e-06 pute = -5.107561938e-13
+ ua1 = 1.732232133e-09 lua1 = 3.603584080e-17 wua1 = 1.030148431e-14 pua1 = -3.605228107e-21
+ ub1 = -4.797891031e-19 lub1 = -3.550784255e-26 wub1 = -1.567823916e-23 pub1 = 3.552404194e-30
+ uc1 = -6.033673320e-11 luc1 = -2.828226037e-18 wuc1 = -1.198373152e-15 puc1 = 2.829516330e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.098241487e+00 lvth0 = 1.801766388e-09 wvth0 = 5.431763791e-07 pvth0 = -1.802588390e-13
+ k1 = 4.964210488e-01 lk1 = -7.181586072e-09 wk1 = -1.572856055e-07 pk1 = 7.184862455e-13
+ k2 = -7.401941116e-03 lk2 = 4.897821019e-09 wk2 = 1.391991276e-06 pk2 = -4.900055503e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.336286821e-01 ldsub = 1.871111750e-08 wdsub = 1.169678066e-05 pdsub = -1.871965389e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.365884236e-01 lvoff = 3.266690915e-09 wvoff = 1.220180774e-06 pvoff = -3.268181244e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.231801296e+00 lnfactor = -6.985855141e-08 wnfactor = -3.574172821e-05 pnfactor = 6.989042228e-12
+ eta0 = -1.428617406e-01 leta0 = 1.975380374e-08 weta0 = 1.434271451e-05 peta0 = -1.976281582e-12
+ etab = -1.435743743e-02 letab = 2.577442070e-09 wetab = 1.386375947e-06 petab = -2.578617951e-13
+ u0 = 1.376773650e-02 lu0 = -4.986372200e-11 wu0 = -9.735121297e-08 pu0 = 4.988647083e-15
+ ua = -6.974822802e-10 lua = -1.670346527e-17 wua = -1.865696578e-14 pua = 1.671108572e-21
+ ub = 1.792656427e-18 lub = 1.640004684e-26 wub = 8.708418478e-24 pub = -1.640752887e-30
+ uc = -7.907655520e-11 luc = 2.977100152e-19 wuc = 6.290253630e-16 puc = -2.978458364e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.028525324e+04 lvsat = 1.046951598e-03 wvsat = 6.703397593e-01 pvsat = -1.047429239e-7
+ a0 = 1.833811615e+00 la0 = 8.735570988e-10 wa0 = -8.221010392e-06 pa0 = -8.739556330e-14
+ ags = 7.648665260e-01 wags = 3.418067077e-6
+ a1 = 0.0
+ a2 = 8.290347267e-01 la2 = -4.334781278e-09 wa2 = -2.904797287e-06 pa2 = 4.336758892e-13
+ b0 = 8.294764088e-25 lb0 = -1.541747801e-31 wb0 = -8.298548325e-29 pb0 = 1.542451177e-35
+ b1 = 0.0
+ keta = -2.919241805e-02 lketa = -4.866751944e-09 wketa = -2.850935756e-06 pketa = 4.868972254e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.722944029e-01 lpclm = 5.512430626e-09 wpclm = 3.680490053e-06 ppclm = -5.514945507e-13
+ pdiblc1 = 2.985345433e-01 lpdiblc1 = 1.675311901e-08 wpdiblc1 = 9.150718511e-06 ppdiblc1 = -1.676076212e-12
+ pdiblc2 = -2.508230397e-03 lpdiblc2 = 3.863098635e-10 wpdiblc2 = 2.753350487e-07 ppdiblc2 = -3.864861058e-14
+ pdiblcb = 1.424476603e-02 lpdiblcb = -4.858170014e-10 wpdiblcb = -1.579175176e-06 ppdiblcb = 4.860386408e-14
+ drout = 7.214186447e-01 ldrout = -3.035611431e-08 wdrout = -1.614922871e-05 pdrout = 3.036996337e-12
+ pscbe1 = 8.000479988e+08 lpscbe1 = -7.481570262e-03 wpscbe1 = -4.802068072e+00 ppscbe1 = 7.484983504e-7
+ pscbe2 = 8.717893628e-09 lpscbe2 = -1.702259894e-17 wpscbe2 = -4.541363702e-15 ppscbe2 = 1.703036499e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -4.486325314e-09 lalpha0 = 6.495211042e-16 walpha0 = 4.588417687e-13 palpha0 = -6.498174287e-20
+ alpha1 = 1.075759376e-10 walpha1 = -7.579393929e-16
+ beta0 = 5.698187331e+00 lbeta0 = 1.710045819e-07 wbeta0 = 1.594468366e-04 pbeta0 = -1.710825976e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056778795e-10 wagidl = -4.000419274e-17
+ bgidl = 9.254056573e+08 lbgidl = 8.270917627e+00 wbgidl = 7.462837410e+03 pbgidl = -8.274690985e-4
+ cgidl = 4.177955700e+02 lcgidl = -1.836079550e-05 wcgidl = -1.178493107e-02 pcgidl = 1.836917206e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.283482011e-01 lkt1 = 7.938102615e-10 wkt1 = -2.322858121e-07 pkt1 = -7.941724136e-14
+ kt2 = -3.805906314e-02 lkt2 = -9.151132489e-10 wkt2 = -5.637507627e-07 pkt2 = 9.155307419e-14
+ at = 9.204209485e+04 lat = 6.026373386e-04 wat = -1.142615893e-01 pat = -6.029122738e-8
+ ute = -2.110909566e-01 lute = 8.271722411e-09 wute = 4.449824834e-06 pute = -8.275496137e-13
+ ua1 = 1.959513039e-09 lua1 = -2.581163689e-18 wua1 = -1.243697535e-14 pua1 = 2.582341267e-22
+ ub1 = -7.341682892e-19 lub1 = 8.199072311e-27 wub1 = 9.771284743e-24 pub1 = -8.202812892e-31
+ uc1 = -8.780780837e-11 luc1 = 1.993107584e-18 wuc1 = 1.549987650e-15 puc1 = -1.994016880e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.102819224e+00 lvth0 = -6.819016693e-07 wvth0 = -4.804956195e-08 pvth0 = 4.804421403e-12
+ k1 = 4.350633756e-01 lk1 = 1.508276488e-07 wk1 = 1.062792890e-08 pk1 = -1.062674601e-12
+ k2 = 3.028188102e-02 lk2 = -2.494815317e-07 wk2 = -1.757948228e-08 pk2 = 1.757752569e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.323275629e-01 lvoff = 9.606613573e-07 wvoff = 6.769210207e-08 pvoff = -6.768456794e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.829534605e+00 lnfactor = 4.201762240e-05 wnfactor = 2.960732377e-06 pnfactor = -2.960402848e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.619232567e-02 lu0 = 3.414892212e-07 wu0 = 2.406271788e-08 pu0 = -2.406003970e-12
+ ua = -4.980122662e-10 lua = 2.215036401e-14 wua = 1.560804637e-15 pua = -1.560630920e-19
+ ub = 2.018945184e-18 lub = 3.248703844e-23 wub = 2.289168712e-24 pub = -2.288913927e-28
+ uc = -7.885964217e-11 luc = 1.188813844e-16 wuc = 8.376865321e-18 puc = -8.375932976e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.749829144e+05 lvsat = 2.501430123e+00 wvsat = 1.762609289e-01 pvsat = -1.762413111e-5
+ a0 = 1.577326108e+00 la0 = -7.557599587e-06 wa0 = -5.325391708e-07 pa0 = 5.324798992e-11
+ ags = 4.450855028e-01 lags = -6.263482074e-06 wags = -4.413503932e-07 pags = 4.413012709e-11
+ a1 = 0.0
+ a2 = 8.739259507e-01 la2 = 1.260500183e-05 wa2 = 8.881996389e-07 pa2 = -8.881007823e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.644330552e-02 lketa = 2.327163310e-06 wketa = 1.639813812e-07 pketa = -1.639631301e-11
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.385060400e-01 lpclm = -6.300936432e-06 wpclm = -4.439895795e-07 ppclm = 4.439401635e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.445818285e-03 lpdiblc2 = 2.181538282e-07 wpdiblc2 = 1.537200502e-08 ppdiblc2 = -1.537029412e-12
+ pdiblcb = -1.967595829e-03 lpdiblcb = 1.871643453e-07 wpdiblcb = 1.318836015e-08 ppdiblcb = -1.318689229e-12
+ drout = 0.56
+ pscbe1 = 7.289941771e+08 lpscbe1 = 1.747900731e+03 wpscbe1 = 1.231641866e+02 ppscbe1 = -1.231504784e-2
+ pscbe2 = 9.567980904e-09 lpscbe2 = -6.298139368e-15 wpscbe2 = -4.437924870e-16 ppscbe2 = 4.437430929e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.360966458e-10 lalpha0 = -2.360703682e-14 walpha0 = -1.663447722e-15 palpha0 = 1.663262580e-19
+ alpha1 = 3.713834012e-11 lalpha1 = 6.285466338e-15 walpha1 = 4.428994938e-16 palpha1 = -4.428501991e-20
+ beta0 = 3.797941871e+00 lbeta0 = 9.943365472e-05 wbeta0 = 7.006499276e-06 pbeta0 = -7.005719452e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.341006471e+09 lbgidl = -1.865411064e+04 wbgidl = -1.314444421e+03 pbgidl = 1.314298123e-1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.353864824e-01 lkt1 = -6.302816058e-07 wkt1 = -4.441220256e-08 pkt1 = 4.440725948e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.322217128e-01 lute = 3.155820000e-06 wute = 2.223718982e-07 pute = -2.223471482e-11
+ ua1 = 2.2116e-9
+ ub1 = -8.736257635e-19 lub1 = 8.002685548e-24 wub1 = 5.639017359e-25 pub1 = -5.638389736e-29
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.136933292e+00 wvth0 = 1.923052657e-7
+ k1 = 4.426089572e-01 wk1 = -4.253538653e-8
+ k2 = 1.780085875e-02 wk2 = 7.035708285e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.842677498e-01 wvoff = -2.709191748e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.931585517e+00 wnfactor = -1.184952377e-5
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.327629396e-02 wu0 = -9.630446494e-8
+ ua = 6.101226114e-10 wua = -6.246694835e-15
+ ub = 3.644201561e-18 wub = -9.161773375e-24
+ uc = -7.291226324e-11 wuc = -3.352611857e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.001240616e+05 wvsat = -7.054362909e-1
+ a0 = 1.199235722e+00 wa0 = 2.131342775e-6
+ ags = 1.317370207e-01 wags = 1.766384566e-6
+ a1 = 0.0
+ a2 = 1.504526972e+00 wa2 = -3.554776789e-6
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.997964934e-02 wketa = -6.562907508e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.767162027e-01 wpclm = 1.776947189e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.235958321e-02 wpdiblc2 = -6.152225722e-8
+ pdiblcb = 7.395832182e-03 wpdiblcb = -5.278281424e-8
+ drout = 0.56
+ pscbe1 = 8.164378760e+08 wpscbe1 = -4.929310625e+2
+ pscbe2 = 9.252898593e-09 wpscbe2 = 1.776158380e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.449124269e-10 walpha0 = 6.657495783e-15
+ alpha1 = 3.515866475e-10 walpha1 = -1.772584419e-15
+ beta0 = 8.772392889e+00 wbeta0 = -2.804160225e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 4.077815992e+08 wbgidl = 5.260705265e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.669181100e-01 wkt1 = 1.777477268e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -1.743428532e-01 wute = -8.899828683e-7
+ ua1 = 2.2116e-9
+ ub1 = -4.732686873e-19 wub1 = -2.256862888e-24
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.159218364e+00 lvth0 = 1.780325398e-07 wvth0 = 2.665158394e-07 pvth0 = -5.928586260e-13
+ k1 = 6.151870697e-01 lk1 = -1.378704106e-06 wk1 = -1.210094400e-06 pk1 = 9.327477176e-12
+ k2 = -5.761121188e-02 lk2 = 6.024572286e-07 wk2 = 5.640866218e-07 pk2 = -3.944341102e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.664452026e-01 lvoff = -1.423820120e-07 wvoff = -3.210364377e-07 pvoff = 4.003802980e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 5.558032831e+00 lnfactor = -1.299347616e-05 wnfactor = -1.881212120e-05 pnfactor = 5.562328575e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.403527535e-02 lu0 = -8.595210369e-08 wu0 = -1.458290766e-07 pu0 = 3.956456845e-13
+ ua = 1.689467794e-09 lua = -8.622748347e-15 wua = -1.146320274e-14 pua = 4.167400354e-20
+ ub = 4.242766131e-18 lub = -4.781854536e-24 wub = -1.157016041e-23 pub = 1.924029091e-29
+ uc = -1.289764046e-10 luc = 4.478891366e-16 wuc = 3.105199470e-16 puc = -2.748539291e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.978419404e+05 lvsat = -7.806554309e-01 wvsat = -8.720088870e-01 pvsat = 1.330726816e-6
+ a0 = 5.406787663e-01 la0 = 5.261125905e-06 wa0 = 4.636363967e-06 pa0 = -2.001228865e-11
+ ags = -3.997935880e-01 lags = 4.246328934e-06 wags = 3.747499350e-06 pags = -1.582686846e-11
+ a1 = 0.0
+ a2 = 2.207093597e+00 la2 = -5.612713438e-06 wa2 = -7.099662412e-06 pa2 = 2.831963040e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.245044653e-01 lketa = -1.154589967e-06 wketa = -1.377977688e-06 pketa = 5.765463121e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -9.839923918e-01 lpclm = 6.449224529e-06 wpclm = 3.548950023e-06 ppclm = -1.415630028e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.354622109e-02 lpdiblc2 = -8.936859575e-08 wpdiblc2 = -1.182104019e-07 ppdiblc2 = 4.528742185e-13
+ pdiblcb = 9.804416972e-03 lpdiblcb = -1.924187077e-08 wpdiblcb = -6.500789127e-08 ppdiblcb = 9.766455109e-14
+ drout = 0.56
+ pscbe1 = 6.416216750e+08 lpscbe1 = 1.396583904e+03 wpscbe1 = 3.626911329e+02 ppscbe1 = -6.835454488e-3
+ pscbe2 = 9.812222954e-09 lpscbe2 = -4.468369613e-15 wpscbe2 = 1.730604322e-15 ppscbe2 = 3.639254470e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.787195635e-09 lalpha0 = 7.527778052e-15 walpha0 = 1.329646708e-14 palpha0 = -5.303787866e-20
+ alpha1 = 6.024732552e-10 lalpha1 = -2.004300493e-15 walpha1 = -3.540236621e-15 palpha1 = 1.412154365e-20
+ beta0 = 1.385922935e+01 lbeta0 = -4.063807519e-05 wbeta0 = -6.756341667e-05 pbeta0 = 3.157346375e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.360692841e-09 lagidl = -7.398247122e-14 wagidl = -6.556589074e-14 pagidl = 5.237973775e-19
+ bgidl = 2.400996867e+09 lbgidl = -1.592353766e+04 wbgidl = -7.697605605e+03 pbgidl = 1.035222610e-1
+ cgidl = 300.0
+ egidl = 6.277691851e-01 legidl = -4.216279410e-06 wegidl = -3.718462182e-06 pegidl = 2.970631097e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.390203810e-01 lkt1 = -2.228713302e-07 wkt1 = 5.686108277e-08 pkt1 = 9.657476841e-13
+ kt2 = -4.616153859e-02 lkt2 = 6.551303671e-08 wkt2 = 7.453494696e-08 pkt2 = -5.954500017e-13
+ at = -4.616340251e+05 lat = 3.687934214e+00 wat = 1.408098974e+00 pat = -1.124911965e-5
+ ute = -2.299268933e+00 lute = 1.697575821e-05 wute = 1.406451037e-05 pute = -1.194695024e-10
+ ua1 = -4.928623343e-09 lua1 = 5.704231605e-14 wua1 = 4.885433424e-14 pua1 = -3.902909252e-19
+ ub1 = 4.325482046e-18 lub1 = -3.833659577e-23 wub1 = -3.484290359e-23 pub1 = 2.603256430e-28
+ uc1 = -8.907706144e-11 luc1 = 1.669091133e-15 wuc1 = 1.352086981e-15 puc1 = -1.080164712e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.115092774e+00 lvth0 = 2.021297172e-09 wvth0 = 8.613294943e-08 pvth0 = 1.266652722e-13
+ k1 = 1.423484992e-01 lk1 = 5.073874829e-07 wk1 = 1.567950669e-06 pk1 = -1.753783457e-12
+ k2 = 1.499335278e-01 lk2 = -2.254117573e-07 wk2 = -6.363463596e-07 pk2 = 8.440300048e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.293770610e+00 ldsub = -2.926915574e-06 wdsub = -3.702329134e-06 pdsub = 1.476810961e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.254349972e-01 lvoff = 9.292060973e-08 wvoff = -1.200608205e-07 pvoff = -4.012853123e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.240901309e+00 lnfactor = 4.227000257e-06 wnfactor = 7.434294489e-07 pnfactor = -2.238126358e-11
+ eta0 = 3.585049213e-01 leta0 = -1.110919925e-06 weta0 = -1.405230558e-06 peta0 = 5.605282015e-12
+ etab = -3.134728557e-01 letab = 9.711815699e-07 wetab = 1.228471997e-06 petab = -4.900215095e-12
+ u0 = 2.592742399e-02 lu0 = -1.372223862e-08 wu0 = -4.935111365e-08 pu0 = 1.080763239e-14
+ ua = -5.138352943e-10 lua = 1.659412420e-16 wua = 1.152263293e-15 pua = -8.647450472e-21
+ ub = 3.707973304e-18 lub = -2.648635473e-24 wub = -9.976797850e-24 pub = 1.288457481e-29
+ uc = 7.129056065e-11 luc = -3.509497529e-16 wuc = -9.818053309e-16 puc = 2.406378240e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.928848552e+05 lvsat = -3.619952623e-01 wvsat = -6.962348514e-01 pvsat = 6.295870386e-7
+ a0 = 1.809673839e+00 la0 = 1.992695294e-07 wa0 = 3.493871911e-07 pa0 = -2.912095596e-12
+ ags = 6.035624379e-01 lags = 2.440721825e-07 wags = -9.490079668e-07 pags = 2.906888677e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.730298644e-02 lketa = 8.916942351e-08 wketa = 2.410822573e-07 pketa = -6.927565222e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.735829217e-01 lpclm = 1.432920088e-06 wpclm = 2.697257863e-06 ppclm = -1.075901097e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.962187643e-03 lpdiblc2 = -3.272692266e-09 wpdiblc2 = -8.815648409e-09 ppdiblc2 = 1.651276809e-14
+ pdiblcb = 1.145869460e-02 lpdiblcb = -2.584056916e-08 wpdiblcb = -8.078046494e-08 ppdiblcb = 1.605792971e-13
+ drout = 0.56
+ pscbe1 = 1.181086351e+09 lpscbe1 = -7.552705583e+02 wpscbe1 = -2.684990378e+03 ppscbe1 = 5.321350861e-3
+ pscbe2 = 9.692068049e-09 lpscbe2 = -3.989087317e-15 wpscbe2 = -3.275750079e-15 ppscbe2 = 2.033362233e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.780816322e-03 lalpha0 = -1.109231440e-08 walpha0 = -1.959257995e-08 palpha0 = 7.815225438e-14
+ alpha1 = -1.508771557e-10 lalpha1 = 1.000716360e-15 walpha1 = 1.767585607e-15 palpha1 = -7.050669202e-21
+ beta0 = 6.776916852e+01 lbeta0 = -2.556778142e-04 wbeta0 = -4.538596138e-04 pbeta0 = 1.856619949e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.843987568e-08 lagidl = 3.691038253e-14 wagidl = 1.312250750e-13 pagidl = -2.611762019e-19
+ bgidl = -3.329181833e+09 lbgidl = 6.933400255e+03 wbgidl = 3.050177876e+04 pbgidl = -4.885011737e-2
+ cgidl = 300.0
+ egidl = -9.555383702e-01 legidl = 2.099328598e-06 wegidl = 7.436924363e-06 pegidl = -1.479107576e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.882472553e-01 lkt1 = 3.723752719e-07 wkt1 = 8.040359317e-07 pkt1 = -2.014635656e-12
+ kt2 = -2.943788167e-02 lkt2 = -1.195456665e-09 wkt2 = -5.339700739e-08 pkt2 = -8.514606699e-14
+ at = 7.379216042e+05 lat = -1.096937249e+00 wat = -2.147199903e+00 pat = 2.932505380e-6
+ ute = 4.316411536e+00 lute = -9.413331140e-06 wute = -3.343546404e-05 pute = 7.000172055e-11
+ ua1 = 1.787229139e-08 lua1 = -3.390756870e-14 wua1 = -1.047961370e-13 pua1 = 2.226008302e-19
+ ub1 = -1.147124632e-17 lub1 = 2.467450012e-23 wub1 = 7.168180679e-23 pub1 = -1.645875785e-28
+ uc1 = 1.047266131e-09 luc1 = -2.863634138e-15 wuc1 = -4.947967883e-15 puc1 = 1.432845273e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.151831237e+00 lvth0 = 7.508932502e-08 wvth0 = 2.669492132e-07 pvth0 = -2.329547703e-13
+ k1 = 3.426293699e-01 lk1 = 1.090548675e-07 wk1 = 1.422595963e-06 pk1 = -1.464691844e-12
+ k2 = 4.309155025e-02 lk2 = -1.291695333e-08 wk2 = -3.964417812e-07 pk2 = 3.668909860e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.708461534e+00 ldsub = 3.044133870e-06 wdsub = 9.982070188e-06 pdsub = -1.244838167e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.404586037e-01 lvoff = -7.608639003e-08 wvoff = -5.761974844e-07 pvoff = 5.059112146e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 5.657363919e+00 lnfactor = -4.556769733e-06 wnfactor = -2.493436669e-05 pnfactor = 2.868853483e-11
+ eta0 = -6.146900923e-01 leta0 = 8.246384413e-07 weta0 = 2.806618621e-06 peta0 = -2.771538461e-12
+ etab = -4.063511457e-01 letab = 1.155904414e-06 wetab = 2.862957363e-06 petab = -8.150994004e-12
+ u0 = 2.493592518e-02 lu0 = -1.175027639e-08 wu0 = -7.657358145e-08 pu0 = 6.494958192e-14
+ ua = 1.764193197e-10 lua = -1.206885452e-15 wua = -8.093219902e-15 pua = 9.740613691e-21
+ ub = 2.635229046e-18 lub = -5.150866001e-25 wub = -2.792691989e-24 pub = -1.403677816e-30
+ uc = -1.277722590e-10 luc = 4.496031725e-17 wuc = 3.259101763e-16 puc = -1.944979013e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.273593820e+04 lvsat = 3.607491425e-02 wvsat = -4.731944871e-01 pvsat = 1.859887492e-7
+ a0 = 6.280821975e-01 la0 = 2.549301697e-06 wa0 = 7.730529304e-06 pa0 = -1.759222771e-11
+ ags = -4.175703062e-01 lags = 2.274972463e-06 wags = 7.721830343e-06 pags = -1.433828151e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.766171263e-02 lketa = -1.394804175e-07 wketa = -7.111568984e-07 pketa = 1.201123367e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.689760276e-01 lpclm = 4.987360150e-08 wpclm = -3.322450308e-06 ppclm = 1.213406018e-12
+ pdiblc1 = 5.326869814e-01 lpdiblc1 = -2.837858568e-07 wpdiblc1 = -6.886815378e-07 ppdiblc1 = 1.369698050e-12
+ pdiblc2 = 2.046297715e-04 lpdiblc2 = 2.228618578e-10 wpdiblc2 = -1.020410556e-09 ppdiblc2 = 1.009053386e-15
+ pdiblcb = -6.075014542e-02 lpdiblcb = 1.177734265e-07 wpdiblcb = 4.157835738e-07 ppdiblcb = -8.270220226e-13
+ drout = -9.238901618e-02 ldrout = 1.297516943e-06 wdrout = 2.580118768e-06 pdrout = -5.131520814e-12
+ pscbe1 = 8.026606526e+08 lpscbe1 = -2.631039524e+00 wpscbe1 = -1.874595240e+01 ppscbe1 = 1.853730995e-5
+ pscbe2 = 6.547310944e-09 lpscbe2 = 2.265425748e-15 wpscbe2 = 1.196539533e-14 ppscbe2 = -9.979034533e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.526342102e-03 lalpha0 = 5.429543773e-09 walpha0 = 3.893651820e-08 palpha0 = -3.825451305e-14
+ alpha1 = 3.522811000e-10 walpha1 = -1.777477268e-15
+ beta0 = -8.153451963e+01 lbeta0 = 4.126781201e-05 wbeta0 = 6.152475333e-04 pbeta0 = -2.696951824e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.369799885e-10 lagidl = -3.656840127e-17 wagidl = -1.865870437e-16 pagidl = 1.845103299e-22
+ bgidl = -1.206890748e+08 lbgidl = 5.521252629e+02 wbgidl = 7.014341783e+03 pbgidl = -2.136658580e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.551411609e-01 lkt1 = -9.124244614e-08 wkt1 = -2.520107908e-07 pkt1 = 8.570398938e-14
+ kt2 = -1.154294599e-02 lkt2 = -3.678615740e-08 wkt2 = -2.021935746e-07 pkt2 = 2.107909617e-13
+ at = 1.326236721e+05 lat = 1.069216493e-01 wat = -6.807401875e-01 pat = 1.590764569e-8
+ ute = 5.080731928e-01 lute = -1.839041260e-06 wute = 3.913726864e-06 pute = -4.280964767e-12
+ ua1 = 2.914363291e-09 lua1 = -4.158194237e-15 wua1 = 9.676223884e-15 pua1 = -5.069814264e-21
+ ub1 = 6.859052361e-23 lub1 = 1.859546029e-24 wub1 = -1.424483372e-23 pub1 = 6.309338986e-30
+ uc1 = -6.961398448e-10 luc1 = 6.037737057e-16 wuc1 = 3.893070716e-15 puc1 = -3.255223712e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.071334021e+00 lvth0 = -4.511956697e-09 wvth0 = -1.584247455e-07 pvth0 = 1.876847762e-13
+ k1 = 4.367941770e-01 lk1 = 1.593811473e-08 wk1 = -1.847848047e-07 pk1 = 1.247987759e-13
+ k2 = 4.316230198e-02 lk2 = -1.298691759e-08 wk2 = -4.659581481e-08 pk2 = 2.093880519e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.731635027e+00 ldsub = -3.576744154e-07 wdsub = -5.154823839e-06 pdsub = 2.520038730e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.511711911e-01 lvoff = 3.339396635e-08 wvoff = 1.697145725e-07 pvoff = -2.316988412e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -2.119297491e+00 lnfactor = 3.133337435e-06 wnfactor = 2.053452112e-05 pnfactor = -1.627428426e-11
+ eta0 = 5.200509789e-01 leta0 = -2.974729618e-07 weta0 = -6.992748246e-07 peta0 = 6.953343906e-13
+ etab = 1.511287979e+00 letab = -7.403913865e-07 wetab = -1.065500945e-05 petab = 5.216517842e-12
+ u0 = 1.280510454e-02 lu0 = 2.455282151e-10 wu0 = 9.133953404e-09 pu0 = -1.980402808e-14
+ ua = -1.736210452e-09 lua = 6.844567498e-16 wua = 7.704838107e-15 pua = -5.881611933e-21
+ ub = 3.124040065e-18 lub = -9.984571528e-25 wub = -9.132687820e-24 pub = 4.865753860e-30
+ uc = -1.379956254e-10 luc = 5.506989761e-17 wuc = 1.835153721e-16 puc = -5.368795118e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.824693803e+05 lvsat = -1.515467946e-01 wvsat = -1.052945333e+00 pvsat = 7.592869684e-7
+ a0 = 5.737345141e+00 la0 = -2.503095150e-06 wa0 = -2.311061305e-05 pa0 = 1.290565273e-11
+ ags = 3.218613641e+00 lags = -1.320740756e-06 wags = -1.628537714e-05 pags = 9.401725753e-12
+ a1 = 0.0
+ a2 = 1.883321980e-01 la2 = 6.048599394e-07 wa2 = 2.931891719e-06 pa2 = -2.899259765e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.978374128e-01 lketa = 8.350890261e-08 wketa = 1.021553884e-06 pketa = -5.123023442e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.098471692e-01 lpclm = 5.038923557e-07 wpclm = 3.434340253e-07 ppclm = -2.411677023e-12
+ pdiblc1 = 1.271271525e+00 lpdiblc1 = -1.014149954e-06 wpdiblc1 = -4.540081969e-06 ppdiblc1 = 5.178232394e-12
+ pdiblc2 = 2.136751842e-03 lpdiblc2 = -1.687755694e-09 wpdiblc2 = -1.441310473e-08 ppdiblc2 = 1.425268687e-14
+ pdiblcb = 1.398423604e-01 lpdiblcb = -8.058648472e-08 wpdiblcb = -8.317322400e-07 ppdiblcb = 4.066089402e-13
+ drout = 8.712825320e-01 ldrout = 3.445710587e-07 wdrout = -8.693426349e-07 pdrout = -1.720451917e-12
+ pscbe1 = 9.413387817e+08 lpscbe1 = -1.397656810e+02 wpscbe1 = -7.131420662e+02 ppscbe1 = 7.052047950e-4
+ pscbe2 = 8.935615814e-09 lpscbe2 = -9.629728971e-17 wpscbe2 = 9.730156006e-16 ppscbe2 = 8.910000061e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.058038197e-05 lalpha0 = 3.450468022e-11 walpha0 = 4.972833965e-10 palpha0 = -2.431069341e-16
+ alpha1 = 5.989464227e-10 lalpha1 = -2.439199377e-16 walpha1 = -3.515387893e-15 palpha1 = 1.718567679e-21
+ beta0 = -8.738881919e+01 lbeta0 = 4.705695321e-05 wbeta0 = 6.760164052e-04 pbeta0 = -3.297876966e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -2.886618402e+08 lbgidl = 7.182284913e+02 wbgidl = 9.677666015e+03 pbgidl = -4.770340014e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.077320673e-01 lkt1 = -3.923687649e-08 wkt1 = -3.105783279e-07 pkt1 = 1.436196698e-13
+ kt2 = -6.831870466e-02 lkt2 = 1.935768709e-08 wkt2 = 4.885926778e-08 pkt2 = -3.746766260e-14
+ at = 4.632962301e+05 lat = -2.200705231e-01 wat = -1.499581909e+00 pat = 8.256356592e-7
+ ute = -2.565694443e+00 lute = 1.200515342e-06 wute = -8.215953660e-07 pute = 4.016533266e-13
+ ua1 = -5.201764567e-09 lua1 = 3.867601118e-15 wua1 = 9.982821821e-15 pua1 = -5.372999766e-21
+ ub1 = 6.150217945e-18 lub1 = -4.222152163e-24 wub1 = -1.832412900e-23 pub1 = 1.034323171e-29
+ uc1 = 5.474096425e-11 luc1 = -1.387498000e-16 wuc1 = 9.565556876e-16 puc1 = -3.513920959e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.076884406e+00 lvth0 = -1.798540392e-09 wvth0 = 2.736659916e-07 pvth0 = -2.355142242e-14
+ k1 = 2.357404101e-01 lk1 = 1.142272698e-07 wk1 = -8.598265993e-08 pk1 = 7.649737133e-14
+ k2 = 9.900206785e-02 lk2 = -4.028530393e-08 wk2 = 2.648302626e-08 pk2 = -1.478724785e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.394750045e+00 ldsub = -1.929814546e-07 wdsub = -6.507213452e-07 pdsub = 3.181181441e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -9.187540177e-02 lvoff = -4.448096620e-08 wvoff = -7.150583500e-07 pvoff = 2.008400974e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 5.491772705e+00 lnfactor = -5.874864520e-07 wnfactor = -1.902762705e-05 pnfactor = 3.066463115e-12
+ eta0 = -6.411277589e-01 leta0 = 2.701924878e-07 weta0 = 1.413919628e-06 peta0 = -3.377429816e-13
+ etab = -5.674954363e-03 letab = 1.206282599e-09 wetab = 3.041347972e-08 petab = -7.264867901e-15
+ u0 = 2.099426325e-02 lu0 = -3.757905802e-09 wu0 = -6.178232228e-08 pu0 = 1.486481162e-14
+ ua = 1.245578941e-09 lua = -7.732506304e-16 wua = -9.535092306e-15 pua = 2.546472848e-21
+ ub = 2.762732061e-19 lub = 3.937306315e-25 wub = 2.510336035e-24 pub = -8.261712118e-31
+ uc = -8.230069429e-11 luc = 2.784231663e-17 wuc = 3.745930698e-16 puc = -1.471001053e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.333785337e+05 lvsat = 5.174877511e-02 wvsat = 1.068129581e+00 pvsat = -2.776429249e-7
+ a0 = 3.687733935e-01 la0 = 1.214385206e-07 wa0 = 7.071224328e-06 pa0 = -1.849342110e-12
+ ags = -2.019838439e+00 lags = 1.240181312e-06 wags = 1.158989026e-05 pags = -4.225656222e-12
+ a1 = 0.0
+ a2 = 2.023335604e+00 la2 = -2.922181757e-07 wa2 = -5.863783439e-06 pa2 = 1.400681950e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.775409284e-04 lketa = -1.307219194e-08 wketa = 1.671825008e-07 pketa = -9.462580599e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.119052267e+00 lpclm = -2.827997406e-07 wpclm = -7.541388585e-06 ppclm = 1.442976206e-12
+ pdiblc1 = -2.057828753e+00 lpdiblc1 = 6.133472987e-07 wpdiblc1 = 1.274411926e-05 ppdiblc1 = -3.271495060e-12
+ pdiblc2 = -1.052193208e-02 lpdiblc2 = 4.500695113e-09 wpdiblc2 = 2.780959603e-08 ppdiblc2 = -6.388724848e-15
+ pdiblcb = -0.025
+ drout = 2.260665214e+00 ldrout = -3.346564528e-07 wdrout = -6.578929859e-06 pdrout = 1.070793990e-12
+ pscbe1 = 5.173224367e+08 lpscbe1 = 6.752318955e+01 wpscbe1 = 1.426284132e+03 ppscbe1 = -3.406964907e-4
+ pscbe2 = 1.613274885e-08 lpscbe2 = -3.614759719e-15 wpscbe2 = 5.466712571e-15 ppscbe2 = -1.305833632e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.268145045e-08 lalpha0 = 2.580326768e-14 walpha0 = 2.663152476e-13 palpha0 = -1.301935351e-19
+ alpha1 = 4.365975454e-10 lalpha1 = -1.645524420e-16 walpha1 = -1.698343980e-15 palpha1 = 8.302694217e-22
+ beta0 = -1.744304970e+01 lbeta0 = 1.286256489e-05 wbeta0 = 1.357789499e-04 pbeta0 = -6.568181191e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.015572358e+09 lbgidl = 8.062751900e+01 wbgidl = 5.891334639e+02 pbgidl = -3.272291055e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.325448675e-01 lkt1 = -2.710664286e-08 wkt1 = -3.636361277e-07 pkt1 = 1.695580364e-13
+ kt2 = -2.386568597e-02 lkt2 = -2.374060162e-09 wkt2 = -2.358096856e-08 pkt2 = -2.053804258e-15
+ at = -3.680751891e+04 lat = 2.441519666e-02 wat = 5.055652706e-01 pat = -1.546206427e-7
+ ute = -1.118874046e-01 lute = 9.226954631e-10 wute = -3.906191155e-07 pute = 1.909619670e-13
+ ua1 = 4.214192790e-09 lua1 = -7.355779551e-16 wua1 = -2.430299690e-15 pua1 = 6.954029476e-22
+ ub1 = -4.504795523e-18 lub1 = 9.867642713e-25 wub1 = 8.025112197e-24 pub1 = -2.538121832e-30
+ uc1 = -3.249743350e-10 luc1 = 4.688161836e-17 wuc1 = 9.759192973e-17 puc1 = 6.852951647e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.111672278e-01 lvth0 = -4.138340265e-08 wvth0 = 4.762797134e-07 pvth0 = -7.194976214e-14
+ k1 = -4.824469119e-01 lk1 = 2.857806754e-07 wk1 = 4.636705560e-06 pk1 = -1.051611164e-12
+ k2 = 3.316496711e-01 lk2 = -9.585783692e-08 wk2 = -1.452378614e-06 pk2 = 3.384684322e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.287085407e+00 ldsub = -6.450036024e-07 wdsub = -1.632919047e-05 pdsub = 4.063234064e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.857338210e-01 lvoff = -2.206100561e-08 wvoff = 7.244497016e-08 pvoff = 1.272917935e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.484294219e+00 lnfactor = -1.063440066e-06 wnfactor = -3.698291395e-05 pnfactor = 7.355442497e-12
+ eta0 = 0.49
+ etab = -6.249997450e-04 letab = -6.090131524e-17 wetab = -1.286411089e-15 petab = 3.072850160e-22
+ u0 = 2.032239532e-02 lu0 = -3.597416711e-09 wu0 = -7.448519702e-08 pu0 = 1.789914731e-14
+ ua = 1.888973283e-09 lua = -9.269382369e-16 wua = -2.064889989e-14 pua = 5.201228065e-21
+ ub = -3.001704319e-19 lub = 5.314257234e-25 wub = 1.346828750e-23 pub = -3.443697078e-30
+ uc = 6.421360169e-11 luc = -7.155553250e-18 wuc = -2.659910428e-16 puc = 5.916221718e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.802268818e+05 lvsat = -2.316215048e-02 wvsat = -7.975123405e-01 pvsat = 1.680029609e-7
+ a0 = 3.322190226e+00 la0 = -5.840441581e-07 wa0 = -1.488909283e-05 pa0 = 3.396318850e-12
+ ags = 7.808785771e+00 lags = -1.107582153e-06 wags = -2.081684479e-05 pags = 3.515340579e-12
+ a1 = 0.0
+ a2 = 3.954555545e-02 la2 = 1.816497532e-07 wa2 = 6.639653440e-06 pa2 = -1.586014017e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.147414154e-01 lketa = -8.832077004e-08 wketa = -2.821847028e-06 pketa = 6.193636776e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.187796882e+00 lpclm = -6.035076660e-08 wpclm = -2.958277732e-06 ppclm = 3.482085171e-13
+ pdiblc1 = 8.626234743e-01 lpdiblc1 = -8.426112488e-08 wpdiblc1 = -3.993892463e-06 ppdiblc1 = 7.267138002e-13
+ pdiblc2 = 5.604675091e-03 lpdiblc2 = 6.485324593e-10 wpdiblc2 = 8.874469673e-09 ppdiblc2 = -1.865691216e-15
+ pdiblcb = 7.680222456e-01 lpdiblcb = -1.894292238e-07 wpdiblcb = -3.031142565e-06 ppdiblcb = 7.240490246e-13
+ drout = 5.179002047e-01 ldrout = 8.163782487e-08 wdrout = -7.802466472e-08 pdrout = -4.820772341e-13
+ pscbe1 = 7.987271780e+08 lpscbe1 = 3.040389852e-01 wpscbe1 = 1.070594185e+01 ppscbe1 = -2.557328329e-6
+ pscbe2 = -5.473616084e-08 lpscbe2 = 1.331369674e-14 wpscbe2 = 2.519228739e-13 ppscbe2 = -6.017681689e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.612550594e-08 lalpha0 = -2.576149992e-15 walpha0 = -3.331397454e-13 palpha0 = 1.299827908e-20
+ alpha1 = -2.522811000e-10 walpha1 = 1.777477268e-15
+ beta0 = 4.221536133e+01 lbeta0 = -1.388039759e-06 wbeta0 = -1.722413283e-04 pbeta0 = 7.894991965e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -8.366471076e+08 lbgidl = 5.230671827e+02 wbgidl = 1.201349619e+04 pbgidl = -3.056166629e-3
+ cgidl = 2.432791151e+03 lcgidl = -5.094598222e-04 wcgidl = -1.076125795e-02 pcgidl = 2.570541687e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.317930322e-01 lkt1 = -2.728623376e-08 wkt1 = -1.050357328e-07 pkt1 = 1.077861601e-13
+ kt2 = 1.271108929e-02 lkt2 = -1.111115447e-08 wkt2 = -1.098084317e-07 pkt2 = 1.854334986e-14
+ at = 1.130772970e+05 lat = -1.138778932e-02 wat = -2.692591021e-01 pat = 3.046165526e-8
+ ute = -1.407145244e+00 lute = 3.103209356e-07 wute = 1.154956856e-05 pute = -2.661190664e-12
+ ua1 = 2.961418227e-09 lua1 = -4.363276953e-16 wua1 = 1.641103723e-15 pua1 = -2.771331857e-22
+ ub1 = -1.445563025e-18 lub1 = 2.560054044e-25 wub1 = -8.873761167e-24 pub1 = 1.498512048e-30
+ uc1 = -4.166419301e-10 luc1 = 6.877825681e-17 wuc1 = 1.312018582e-15 puc1 = -2.215605779e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.767872713e-01 lvth0 = -3.335263729e-08 wvth0 = -3.125441138e-07 pvth0 = 6.742580095e-14
+ k1 = 2.065713039e+00 lk1 = -1.590765159e-07 wk1 = -1.121392378e-05 pk1 = 1.788680505e-12
+ k2 = -1.131625526e-01 lk2 = -2.283051622e-08 wk2 = 2.137140567e-06 pk2 = -2.946421674e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.065081894e+00 ldsub = 8.424817669e-07 wdsub = 4.902949247e-05 pdsub = -7.675941999e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.555867589e-01 lvoff = -1.129830281e-08 wvoff = 1.354035863e-06 pvoff = -2.241986842e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -9.829184027e+00 lnfactor = 2.047560524e-06 wnfactor = 4.923541532e-05 pnfactor = -7.929492192e-12
+ eta0 = 1.891873008e+00 leta0 = -2.605661360e-07 weta0 = 6.742604475e-09 peta0 = -1.253247894e-15
+ etab = 3.055636466e-01 letab = -5.691128375e-08 wetab = -8.676670805e-07 petab = 1.612732803e-13
+ u0 = -3.551457769e-02 lu0 = 6.418852566e-09 wu0 = 2.498733440e-07 pu0 = -4.058748271e-14
+ ua = -1.465795725e-08 lua = 2.055325654e-15 wua = 7.970326381e-14 pua = -1.292762537e-20
+ ub = 1.121124418e-17 lub = -1.554702733e-24 wub = -5.765139062e-23 pub = 9.428643424e-30
+ uc = 2.753551710e-10 luc = -4.712078022e-17 wuc = -1.868166604e-15 puc = 3.043081744e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.207709184e+04 lvsat = 1.582577500e-02 wvsat = 1.321089930e+00 pvsat = -2.088689272e-7
+ a0 = -7.273413919e-01 la0 = 1.098470525e-07 wa0 = 9.823905579e-06 pa0 = -8.551816199e-13
+ ags = 1.25
+ a1 = 0.0
+ a2 = 2.924370978e+00 la2 = -3.362662212e-07 wa2 = -1.766774448e-05 pa2 = 2.772339345e-12
+ b0 = -3.857065301e-23 lb0 = 7.169127274e-30 wb0 = 1.946129354e-28 pb0 = -3.617270630e-35
+ b1 = 0.0
+ keta = -1.000116229e+00 lketa = 1.471806431e-07 wketa = 3.989826405e-06 pketa = -5.843712461e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.867697356e+00 lpclm = -1.927993284e-07 wpclm = -5.446429493e-06 ppclm = 8.457351416e-13
+ pdiblc1 = 9.676613367e-01 lpdiblc1 = -1.122670085e-07 wpdiblc1 = 4.436304055e-06 ppdiblc1 = -7.670491633e-13
+ pdiblc2 = 3.218940421e-02 lpdiblc2 = -4.227483929e-09 wpdiblc2 = 3.086863098e-08 ppdiblc2 = -6.141563533e-15
+ pdiblcb = -2.420745796e+00 lpdiblcb = 3.841974125e-07 wpdiblcb = 1.557684790e-05 ppdiblcb = -2.661728760e-12
+ drout = 1.008278222e+00 ldrout = -1.290326457e-09 wdrout = -1.817033286e-05 pdrout = 2.832209783e-12
+ pscbe1 = 8.032688971e+08 lpscbe1 = -5.095229859e-01 wpscbe1 = -2.749529989e+01 ppscbe1 = 4.285692394e-6
+ pscbe2 = 9.832662827e-08 lpscbe2 = -1.379580529e-14 wpscbe2 = -6.358906359e-13 ppscbe2 = 9.878313094e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.133641271e-07 lalpha0 = -3.020273135e-14 walpha0 = -1.076050171e-12 palpha0 = 1.523915657e-19
+ alpha1 = -2.522811000e-10 walpha1 = 1.777477268e-15
+ beta0 = 6.333469369e+01 lbeta0 = -5.453222852e-06 wbeta0 = -2.466382006e-04 pbeta0 = 2.251792078e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 4.621900562e+09 lbgidl = -4.388563421e+02 wbgidl = -1.858126842e+04 pbgidl = 2.322820559e-3
+ cgidl = -5.177494006e+03 lcgidl = 8.537769907e-04 wcgidl = 2.763736426e-02 pcgidl = -4.307835967e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.235353412e-01 lkt1 = 4.278002715e-08 wkt1 = 2.552053396e-06 pkt1 = -3.752362548e-13
+ kt2 = -7.634695936e-01 lkt2 = 1.320389985e-07 wkt2 = 4.547217630e-06 pkt2 = -8.451913409e-13
+ at = 4.123296582e+05 lat = -6.815622480e-02 wat = -2.370886692e+00 pat = 4.241577244e-7
+ ute = 5.016015031e+00 lute = -8.523121187e-07 wute = -3.237838811e-05 pute = 5.235798830e-12
+ ua1 = -2.752956097e-09 lua1 = 5.818783204e-16 wua1 = 2.076530087e-14 pua1 = -3.859646472e-21
+ ub1 = 4.684208350e-18 lub1 = -8.575633536e-25 wub1 = -2.840454891e-23 pub1 = 5.279553506e-30
+ uc1 = 4.806005855e-10 luc1 = -9.106836066e-17 wuc1 = -2.454803035e-15 puc1 = 4.562742401e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108465043e+00 lvth0 = -1.173826690e-07 wvth0 = -1.956289651e-08 pvth0 = 1.956071916e-12
+ k1 = 4.568416918e-01 lk1 = -2.026761573e-06 wk1 = -9.925722216e-08 pk1 = 9.924617483e-12
+ k2 = 1.854189619e-02 lk2 = 9.243862853e-07 wk2 = 4.165604346e-08 pk2 = -4.165140714e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.207646451e-01 lvoff = -1.955017313e-07 wvoff = 9.349989435e-09 pvoff = -9.348948781e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.401997552e+00 lnfactor = -1.522230072e-05 wnfactor = 7.230074105e-08 pnfactor = -7.229269398e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.052377368e-02 lu0 = -9.160737090e-08 wu0 = 2.207868500e-09 pu0 = -2.207622764e-13
+ ua = -1.818148443e-10 lua = -9.465858904e-15 wua = -3.460803100e-17 pua = 3.460417912e-21
+ ub = 2.410868435e-18 lub = -6.700924611e-24 wub = 3.116721315e-25 pub = -3.116374424e-29
+ uc = -8.847927211e-11 luc = 1.080737311e-15 wuc = 5.691388173e-17 puc = -5.690754722e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.099163535e+05 lvsat = -9.915249786e-1
+ a0 = 1.470922768e+00 la0 = 3.081550225e-06 wa0 = 4.331866504e-09 pa0 = -4.331384368e-13
+ ags = 3.569179816e-01 lags = 2.552288740e-06 wags = 3.509591313e-09 pags = -3.509200695e-13
+ a1 = 0.0
+ a2 = 1.049959676e+00 la2 = -4.996411477e-6
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.230853340e-03 lketa = -1.639811003e-06 wketa = -3.619942751e-08 pketa = 3.619539852e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.635223146e-03 lpclm = 6.884677536e-06 wpclm = 2.213807154e-07 ppclm = -2.213560757e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 4.538308903e-03 lpdiblc2 = -9.106081414e-08 wpdiblc2 = -2.315336763e-10 ppdiblc2 = 2.315079066e-14
+ pdiblcb = 1.230263679e-03 lpdiblcb = -1.325860133e-07 wpdiblcb = -2.946830134e-09 ppdiblcb = 2.946502152e-13
+ drout = 0.56
+ pscbe1 = 7.806156748e+08 lpscbe1 = -3.413674501e+03 wpscbe1 = -1.372983783e+02 ppscbe1 = 1.372830970e-2
+ pscbe2 = 9.387039523e-09 lpscbe2 = 1.179398485e-14 wpscbe2 = 4.691693253e-16 ppscbe2 = -4.691171067e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.360966458e-10 lalpha0 = 2.360703682e-14 walpha0 = 7.190611385e-16 palpha0 = -7.189811070e-20
+ alpha1 = 1.628616599e-10 lalpha1 = -6.285466338e-15 walpha1 = -1.914528543e-16 palpha1 = 1.914315456e-20
+ beta0 = 5.104848607e+00 lbeta0 = -3.124247305e-05 wbeta0 = 4.123418947e-07 pbeta0 = -4.122960010e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.174766428e-10 lagidl = -1.747469768e-15 wagidl = -8.818053353e-17 pagidl = 8.817071904e-21
+ bgidl = 9.091179662e+08 lbgidl = 2.452993290e+04 wbgidl = 8.647017195e+02 pbgidl = -8.646054782e-2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.532633165e-01 lkt1 = 1.157202834e-06 wkt1 = 4.578754482e-08 pkt1 = -4.578244866e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -2.801439377e-01 lute = -2.051377888e-06 wute = -4.039286973e-08 pute = 4.038837400e-12
+ ua1 = 2.320991131e-09 lua1 = -1.093789553e-14 wua1 = -5.519462950e-16 pua1 = 5.518848634e-20
+ ub1 = -1.051129558e-18 lub1 = 2.575108939e-23 wub1 = 1.459518787e-24 pub1 = -1.459356343e-28
+ uc1 = 2.362916267e-10 luc1 = -1.164286668e-14 wuc1 = -5.875204336e-16 puc1 = 5.874550426e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.114337444e+00 wvth0 = 7.829515728e-8
+ k1 = 3.554471871e-01 wk1 = 3.972499582e-7
+ k2 = 6.478694583e-02 wk2 = -1.667169518e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.305451745e-01 wvoff = -3.742078241e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.640458719e+00 wnfactor = -2.893639953e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.594085474e-02 wu0 = -8.836391451e-9
+ ua = -6.553713237e-10 wua = 1.385092044e-16
+ ub = 2.075635647e-18 wub = -1.247382695e-24
+ uc = -3.441231829e-11 wuc = -2.277822878e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.625086071e+00 wa0 = -1.733711412e-8
+ ags = 4.846034756e-01 wags = -1.404618195e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.880534994e-02 wketa = 1.448783348e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.510607727e-01 wpclm = -8.860159295e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.726698156e-05 wpdiblc2 = 9.266503862e-10
+ pdiblcb = -5.402728247e-03 wpdiblcb = 1.179388383e-8
+ drout = 0.56
+ pscbe1 = 6.098369114e+08 wpscbe1 = 5.494993096e+2
+ pscbe2 = 9.977067116e-09 wpscbe2 = -1.877722254e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.044912427e-09 walpha0 = -2.877846075e-15
+ alpha1 = -1.515866475e-10 walpha1 = 7.662378286e-16
+ beta0 = 3.541855149e+00 wbeta0 = -1.650285963e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.005450403e-11 wagidl = 3.529185333e-16
+ bgidl = 2.136297537e+09 wbgidl = -3.460732776e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.953709577e-01 wkt1 = -1.832521591e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.827699434e-01 wute = 1.616614435e-7
+ ua1 = 1.773791837e-09 wua1 = 2.209014496e-15
+ ub1 = 2.371418346e-19 wub1 = -5.841325846e-24
+ uc1 = -3.461758503e-10 wuc1 = 2.351390283e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.125470039e+00 lvth0 = 8.893685036e-08 wvth0 = 9.623454736e-08 pvth0 = -1.433154552e-13
+ k1 = 2.581902401e-01 lk1 = 7.769731063e-07 wk1 = 5.911766575e-07 pk1 = -1.549255190e-12
+ k2 = 1.025307909e-01 lk2 = -3.015306720e-07 wk2 = -2.439293908e-07 pk2 = 6.168401374e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.145729767e-01 lvoff = -1.275998122e-07 wvoff = -7.820188227e-08 pvoff = 3.257949053e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.016191491e+00 lnfactor = -3.001680267e-06 wnfactor = -9.413286141e-07 pnfactor = 5.208460584e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.366151088e-02 lu0 = 1.820938180e-08 wu0 = 7.425457624e-09 pu0 = -1.299137982e-13
+ ua = -1.284830365e-09 lua = 5.028666453e-15 wua = 3.543981481e-15 pua = -2.720587530e-20
+ ub = 2.417371494e-18 lub = -2.730083250e-24 wub = -2.359909068e-24 pub = 8.887828571e-30
+ uc = 4.661972086e-11 luc = -6.473544266e-16 wuc = -5.754717266e-16 puc = 2.777645727e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.307415459e+05 lvsat = -5.626484918e-01 wvsat = -2.888346007e-02 pvsat = 2.307462077e-7
+ a0 = 1.131699728e+00 la0 = 3.941599354e-06 wa0 = 1.654295602e-06 pa0 = -1.335445646e-11
+ ags = 1.703447475e-01 lags = 2.510572125e-06 wags = 8.707968212e-07 pags = -7.068895723e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.559908778e-02 lketa = -1.055031116e-07 wketa = 8.577518185e-08 pketa = 4.721674059e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.009301966e-02 lpclm = 2.244614854e-06 wpclm = -1.769566520e-06 ppclm = 7.058570803e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.488876802e-04 lpdiblc2 = 1.850387651e-09 wpdiblc2 = 1.850722368e-09 ppdiblc2 = -7.382290930e-15
+ pdiblcb = -7.090168188e-03 lpdiblcb = 1.348073832e-08 wpdiblcb = 2.023579930e-08 ppdiblcb = -6.744136523e-14
+ drout = 0.56
+ pscbe1 = 6.114112903e+08 lpscbe1 = -1.257750809e+01 wpscbe1 = 5.151213146e+02 ppscbe1 = 2.746413327e-4
+ pscbe2 = 1.168138527e-08 lpscbe2 = -1.361557616e-14 wpscbe2 = -7.700482174e-15 ppscbe2 = 4.651727205e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.987195635e-09 lalpha0 = -7.527778052e-15 walpha0 = -5.747684544e-15 palpha0 = 2.292676645e-20
+ alpha1 = -4.024732552e-10 lalpha1 = 2.004300493e-15 walpha1 = 1.530343600e-15 palpha1 = -6.104341677e-21
+ beta0 = 2.220999188e+00 lbeta0 = 1.055214657e-05 wbeta0 = -8.841306526e-06 pbeta0 = 5.744812845e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.459663969e-09 lagidl = 7.581212722e-14 wagidl = 2.939451563e-14 pagidl = -2.320095438e-19
+ bgidl = 9.867718769e+08 lbgidl = 9.183411057e+03 wbgidl = -5.619608822e+02 pbgidl = -2.315791182e-2
+ cgidl = 300.0
+ egidl = -4.277691851e-01 legidl = 4.216279410e-06 wegidl = 1.607385441e-06 pegidl = -1.284119333e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.022916677e-01 lkt1 = -7.435983468e-07 wkt1 = -6.330203209e-07 pkt1 = 3.593139375e-12
+ kt2 = -3.138933668e-02 lkt2 = -5.250016399e-8
+ at = -1.881185878e+05 lat = 1.502854942e+00 wat = 2.804346631e-02 pat = -2.240356067e-7
+ ute = 9.853518131e-01 lute = -1.092974686e-05 wute = -2.508444332e-06 pute = 2.133112793e-11
+ ua1 = 3.879498199e-09 lua1 = -1.682221438e-14 wua1 = 4.411882410e-15 pua1 = -1.759842539e-20
+ ub1 = -7.594419955e-20 lub1 = 2.501203626e-24 wub1 = -1.263497049e-23 pub1 = 5.427354390e-29
+ uc1 = -7.518597356e-10 luc1 = 3.240955820e-15 wuc1 = 4.696237823e-15 puc1 = -1.873268216e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108526780e+00 lvth0 = 2.135239484e-08 wvth0 = 5.300342784e-08 pvth0 = 2.912786055e-14
+ k1 = 2.328244978e-01 lk1 = 8.781537546e-07 wk1 = 1.111442980e-06 pk1 = -3.624529915e-12
+ k2 = 1.053904391e-01 lk2 = -3.129374366e-07 wk2 = -4.115987710e-07 pk2 = 1.285651498e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.902044650e-01 lvoff = 1.740843627e-07 wvoff = 2.067414313e-07 pvoff = -8.108069299e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.863805798e-01 lnfactor = 1.504988581e-06 wnfactor = 2.532207040e-06 pnfactor = -8.647021582e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.832293334e-02 lu0 = -4.027312641e-08 wu0 = -6.143794835e-08 pu0 = 1.447733760e-13
+ ua = 1.816042345e-09 lua = -7.340311674e-15 wua = -1.060341858e-14 pua = 2.922626438e-20
+ ub = 1.171029543e-18 lub = 2.241412768e-24 wub = 2.823661404e-24 pub = -1.178876018e-29
+ uc = -2.090983595e-10 luc = 3.726717528e-16 wuc = 4.329311734e-16 puc = -1.244742349e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.704228994e+05 lvsat = -3.220452523e-01 wvsat = -7.833811313e-02 pvsat = 4.280143896e-7
+ a0 = 1.749181885e+00 la0 = 1.478543303e-06 wa0 = 6.546067267e-07 pa0 = -9.366827492e-12
+ ags = 6.995207468e-02 lags = 2.911025446e-06 wags = 1.743388221e-06 pags = -1.054954938e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.699411678e-02 lketa = -2.196046222e-07 wketa = -1.275728226e-08 pketa = 8.652005960e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.170973158e-01 lpclm = 6.268582688e-08 wpclm = 9.640140789e-07 ppclm = -3.845326839e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -4.139009881e-02 lpdiblcb = 1.502987026e-07 wpdiblcb = 1.858745697e-07 ppdiblcb = -7.281528875e-13
+ drout = 0.56
+ pscbe1 = 4.189136490e+08 lpscbe1 = 7.552705583e+02 wpscbe1 = 1.160644974e+03 ppscbe1 = -2.300268628e-3
+ pscbe2 = -2.646401887e-09 lpscbe2 = 4.353610419e-14 wpscbe2 = 5.897950528e-14 ppscbe2 = -2.194605295e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.780816122e-03 lalpha0 = 1.109231440e-08 walpha0 = 8.469315062e-09 palpha0 = -3.378299677e-14
+ alpha1 = 3.508771557e-10 lalpha1 = -1.000716360e-15 walpha1 = -7.640769846e-16 palpha1 = 3.047803762e-21
+ beta0 = -6.443688909e+01 lbeta0 = 2.764417974e-04 wbeta0 = 2.132021790e-04 pbeta0 = -8.282544696e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.893993520e-08 lagidl = -3.747018192e-14 wagidl = -5.737932113e-14 pagidl = 1.141200104e-19
+ bgidl = 5.111398910e+09 lbgidl = -7.269189978e+03 wbgidl = -1.208620113e+04 pbgidl = 2.281078437e-2
+ cgidl = 300.0
+ egidl = 1.155538370e+00 legidl = -2.099328598e-06 wegidl = -3.214770882e-06 pegidl = 6.393761365e-12
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.589575541e-01 lkt1 = 2.802085073e-07 wkt1 = 6.562511708e-07 pkt1 = -1.549597000e-12
+ kt2 = -3.978791304e-02 lkt2 = -1.899933468e-08 wkt2 = -1.174661393e-09 pkt2 = 4.685571591e-15
+ at = 3.698768720e+05 lat = -7.229164073e-01 wat = -2.901853053e-01 pat = 1.045337593e-6
+ ute = -3.330248395e+00 lute = 6.284621347e-06 wute = 5.146691534e-06 pute = -9.204213873e-12
+ ua1 = -2.323147812e-09 lua1 = 7.919334216e-15 wua1 = -2.897584698e-15 pua1 = 1.155808868e-20
+ ub1 = 2.073574380e-18 lub1 = -6.072946550e-24 wub1 = 3.339761462e-24 pub1 = -9.447585148e-30
+ uc1 = 2.772151415e-11 luc1 = 1.313075607e-16 wuc1 = 1.962688676e-16 puc1 = -7.828909981e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.111237418e+00 lvth0 = 2.674350079e-08 wvth0 = 6.212814514e-08 pvth0 = 1.097998404e-14
+ k1 = 9.173808884e-01 lk1 = -4.833399140e-07 wk1 = -1.477382943e-06 pk1 = 1.524308298e-12
+ k2 = -1.328242626e-01 lk2 = 1.608406371e-07 wk2 = 4.911629141e-07 pk2 = -5.098241348e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.447643867e-02 ldsub = 9.457545454e-07 wdsub = 9.355829091e-07 pdsub = -1.860752781e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.860738934e-01 lvoff = -3.301780716e-08 wvoff = -3.460399749e-07 pvoff = 2.886034253e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.473685144e+00 lnfactor = 3.369161525e-07 wnfactor = -3.825105023e-06 pnfactor = 3.996845661e-12
+ eta0 = -5.995440838e-02 leta0 = 2.783511242e-07 weta0 = 7.632050099e-09 peta0 = -1.517915548e-14
+ etab = -6.357158270e-01 letab = 1.125135237e-06 wetab = 4.020244845e-06 petab = -7.995744365e-12
+ u0 = 3.922510693e-03 lu0 = 8.256142175e-09 wu0 = 2.945216500e-08 pu0 = -3.599524376e-14
+ ua = -3.309524365e-09 lua = 2.853774189e-15 wua = 9.495534245e-15 pua = -1.074793993e-20
+ ub = 3.498445948e-18 lub = -2.387515897e-24 wub = -7.148158180e-24 pub = 8.043892638e-30
+ uc = 2.554573859e-11 luc = -9.400485470e-17 wuc = -4.476744853e-16 puc = 5.066678276e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.413607529e+04 lvsat = 1.444620556e-01 wvsat = 3.183223954e-01 pvsat = -3.608917959e-7
+ a0 = 3.750625831e+00 la0 = -2.502068519e-06 wa0 = -8.024645549e-06 pa0 = 7.895076982e-12
+ ags = 2.571431665e+00 lags = -2.064092267e-06 wags = -7.359543761e-06 pags = 7.554998950e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.817890151e-01 lketa = 2.672606071e-07 wketa = 8.502145011e-07 pketa = -8.511380948e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.207572630e-01 lpclm = -1.434803323e-07 wpclm = -2.070032248e-06 ppclm = 2.188996880e-12
+ pdiblc1 = 3.769956971e-01 lpdiblc1 = 2.586386786e-08 wpdiblc1 = 9.687783153e-08 ppdiblc1 = -1.926774128e-13
+ pdiblc2 = 2.392950000e-06 lpdiblc2 = 4.228477835e-10
+ pdiblcb = 9.270092676e-02 lpdiblcb = -1.163909154e-07 wpdiblcb = -3.584725320e-07 ppdiblcb = 3.544827327e-13
+ drout = 8.523031487e-01 ldrout = -5.813529634e-07 wdrout = -2.186440802e-06 pdrout = 4.348546518e-12
+ pscbe1 = 7.973393474e+08 lpscbe1 = 2.631039524e+00 wpscbe1 = 8.103342053e+00 ppscbe1 = -8.013151856e-6
+ pscbe2 = 2.928315775e-08 lpscbe2 = -1.996763908e-14 wpscbe2 = -1.027510935e-13 ppscbe2 = 1.022006065e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.526342302e-03 lalpha0 = -5.429543773e-09 walpha0 = -1.683114939e-08 palpha0 = 1.653633796e-14
+ alpha1 = -1.522811000e-10 walpha1 = 7.683528683e-16
+ beta0 = 9.158106374e+01 lbeta0 = -3.385762846e-05 wbeta0 = -2.582282627e-04 pbeta0 = 1.093593929e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.270113134e+09 lbgidl = 3.706280642e+02 wbgidl = -3.120438703e+00 pbgidl = -1.220892321e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.451299616e-01 lkt1 = -1.450667767e-07 wkt1 = -3.025235182e-07 pkt1 = 3.572812157e-13
+ kt2 = -3.823071454e-02 lkt2 = -2.209640007e-08 wkt2 = -6.753718248e-08 pkt2 = 1.366719989e-13
+ at = -1.046632834e+05 lat = 2.208822715e-01 wat = 5.165200953e-01 pat = -5.590945767e-7
+ ute = 3.238636071e+00 lute = -6.780035903e-06 wute = -9.863661269e-06 pute = 2.064942651e-11
+ ua1 = 7.889564179e-09 lua1 = -1.239242228e-14 wua1 = -1.542675917e-14 pua1 = 3.647698791e-20
+ ub1 = -4.796816849e-18 lub1 = 7.591368453e-24 wub1 = 9.958436984e-24 pub1 = -2.261127033e-29
+ uc1 = -4.245343738e-11 luc1 = 2.708764165e-16 wuc1 = 5.948161973e-16 puc1 = -1.575549826e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.131545913e+00 lvth0 = 4.682596217e-08 wvth0 = 1.453816979e-07 pvth0 = -7.134695664e-14
+ k1 = 5.026836058e-01 lk1 = -7.325821210e-08 wk1 = -5.172379558e-07 pk1 = 5.748497248e-13
+ k2 = -7.579439947e-03 lk2 = 3.698978931e-08 wk2 = 2.094278346e-07 pk2 = -2.312247666e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.080841523e+00 ldsub = -3.952099518e-08 wdsub = -1.871165818e-06 pdsub = 9.147568336e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.940924052e-01 lvoff = -2.508854141e-08 wvoff = -1.182834055e-07 pvoff = 6.338178657e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.548172658e+00 lnfactor = -7.256123152e-07 wnfactor = -3.015768944e-06 pnfactor = 3.196517493e-12
+ eta0 = 4.168013260e-01 leta0 = -1.930983189e-07 weta0 = -1.783161045e-07 peta0 = 1.686993961e-13
+ etab = 9.925540395e-01 letab = -4.850119860e-07 wetab = -8.037674077e-06 petab = 3.927969920e-12
+ u0 = 1.907463994e-02 lu0 = -6.727343869e-09 wu0 = -2.249975232e-08 pu0 = 1.537844872e-14
+ ua = 3.717612460e-10 lua = -7.865387138e-16 wua = -2.931190266e-15 pua = 1.540475141e-21
+ ub = 1.347668433e-18 lub = -2.606765365e-25 wub = -1.697880345e-25 pub = 1.143191751e-30
+ uc = -1.585804685e-10 luc = 8.807202769e-17 wuc = 2.873787091e-16 puc = -2.202042248e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.715945267e+04 lvsat = -5.149553097e-03 wvsat = -6.748526583e-02 pvsat = 2.062182600e-8
+ a0 = 1.041351478e+00 la0 = 1.770516104e-07 wa0 = 5.835958862e-07 pa0 = -6.173547263e-13
+ ags = 1.073595718e-01 lags = 3.725547039e-07 wags = -5.871651639e-07 pags = 8.579969271e-13
+ a1 = 0.0
+ a2 = 1.020591357e+00 la2 = -2.181361750e-07 wa2 = -1.267373402e-06 pa2 = 1.253267536e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.316930213e-02 lketa = 1.630631562e-09 wketa = 8.978840231e-08 pketa = -9.917553844e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.388708941e-01 lpclm = -6.250535871e-08 wpclm = -3.075709197e-07 ppclm = 4.461517458e-13
+ pdiblc1 = 1.308749221e+00 lpdiblc1 = -8.955192397e-07 wpdiblc1 = -4.729180260e-06 ppdiblc1 = 4.579666652e-12
+ pdiblc2 = -1.595917611e-03 lpdiblc2 = 2.003369148e-09 wpdiblc2 = 4.420534383e-09 ppdiblc2 = -4.371333835e-15
+ pdiblcb = 1.172588168e-02 lpdiblcb = -3.631712262e-08 wpdiblcb = -1.853049166e-07 ppdiblcb = 1.832424728e-13
+ drout = 2.267188182e-01 ldrout = 3.726861354e-08 wdrout = 2.382882220e-06 pdrout = -1.699199387e-13
+ pscbe1 = 7.869784414e+08 lpscbe1 = 1.287662868e+01 wpscbe1 = 6.570186271e+01 ppscbe1 = -6.497060098e-5
+ pscbe2 = 8.811227077e-09 lpscbe2 = 2.764390048e-16 wpscbe2 = 1.600634151e-15 ppscbe2 = -9.896864416e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.058058197e-05 lalpha0 = -3.450468022e-11 walpha0 = -2.149614687e-10 palpha0 = 1.050882132e-16
+ alpha1 = -3.989464227e-10 lalpha1 = 2.439199377e-16 walpha1 = 1.519602202e-15 palpha1 = -7.428879284e-22
+ beta0 = 1.046580191e+02 lbeta0 = -4.678903733e-05 wbeta0 = -2.929793472e-04 pbeta0 = 1.437236978e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 2.160768431e+09 lbgidl = -5.101142401e+02 wbgidl = -2.681233251e+03 pbgidl = 1.427413095e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.924717974e-01 lkt1 = 6.351445455e-10 wkt1 = 1.169863187e-07 pkt1 = -5.755947671e-14
+ kt2 = -1.062481582e-01 lkt2 = 4.516400942e-08 wkt2 = 2.402369528e-07 pkt2 = -1.676766103e-13
+ at = 1.619462245e+05 lat = -4.275987261e-02 wat = 2.091630816e-02 pat = -6.900685967e-8
+ ute = -6.913338111e+00 lute = 3.258946807e-06 wute = 2.111497117e-05 pute = -9.984413758e-12
+ ua1 = -1.216904515e-08 lua1 = 7.442934724e-15 wua1 = 4.513708600e-14 pua1 = -2.341278166e-20
+ ub1 = 7.951849306e-18 lub1 = -5.015405048e-24 wub1 = -2.741447983e-23 pub1 = 1.434568592e-29
+ uc1 = 8.020344020e-10 luc1 = -5.642122732e-16 wuc1 = -2.814004522e-15 puc1 = 1.795330719e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.010738833e+00 lvth0 = -1.223299500e-08 wvth0 = -6.007956578e-08 pvth0 = 2.909689132e-14
+ k1 = -1.602433399e-01 lk1 = 2.508268838e-07 wk1 = 1.912001661e-06 pk1 = -6.127326464e-13
+ k2 = 2.443993654e-01 lk2 = -8.619508927e-08 wk2 = -7.071367771e-07 pk2 = 2.168561751e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.068204422e+00 ldsub = -3.334309579e-08 wdsub = 9.969044353e-07 pdsub = -4.873566713e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.281271567e-01 lvoff = -8.449972447e-09 wvoff = -2.758349771e-08 pvoff = 1.904132266e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.143836368e+00 lnfactor = -3.907443314e-08 wnfactor = 2.910416189e-06 pnfactor = 2.993833672e-13
+ eta0 = -4.255318186e-01 leta0 = 2.186930855e-07 weta0 = 3.261040085e-07 peta0 = -7.789646451e-14
+ etab = 1.468804215e-03 letab = -5.001470127e-10 wetab = -5.631225722e-09 petab = 1.345130888e-15
+ u0 = 6.814617104e-03 lu0 = -7.337865075e-10 wu0 = 9.762812260e-09 pu0 = -3.937512269e-16
+ ua = -1.740025874e-10 lua = -5.197311486e-16 wua = -2.372420517e-15 pua = 1.267309373e-21
+ ub = -4.313896939e-19 lub = 6.090516102e-25 wub = 6.080935532e-24 pub = -1.912599479e-30
+ uc = 4.643812610e-11 luc = -1.215541264e-17 wuc = -2.749743547e-16 puc = 5.471331752e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.303938881e+04 lvsat = 1.753322526e-03 wvsat = 2.662276988e-02 pvsat = -2.538476941e-8
+ a0 = 2.079580100e+00 la0 = -3.305072156e-07 wa0 = -1.560859625e-06 pa0 = 4.310052396e-13
+ ags = 2.600371964e-01 lags = 2.979151935e-07 wags = 8.649959848e-08 pags = 5.286624347e-13
+ a1 = 0.0
+ a2 = 3.588172864e-01 la2 = 1.053853148e-07 wa2 = 2.534746804e-06 pa2 = -6.054749690e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.248466783e-01 lketa = -6.584124079e-08 wketa = -4.641470125e-07 pketa = 1.716268678e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.911359554e-01 lpclm = 5.860482075e-08 wpclm = 1.177023973e-06 ppclm = -2.796221592e-13
+ pdiblc1 = -1.248307950e+00 lpdiblc1 = 3.545492998e-07 wpdiblc1 = 8.659583286e-06 ppdiblc1 = -1.965698183e-12
+ pdiblc2 = -4.006168681e-03 lpdiblc2 = 3.181668589e-09 wpdiblc2 = -5.066483103e-09 ppdiblc2 = 2.665844032e-16
+ pdiblcb = -9.845176336e-02 lpdiblcb = 1.754542271e-08 wpdiblcb = 3.706098331e-07 ppdiblcb = -8.852757084e-14
+ drout = 1.595081483e-01 ldrout = 7.012589376e-08 wdrout = 4.022714455e-06 pdrout = -9.715847233e-13
+ pscbe1 = 8.258287353e+08 lpscbe1 = -6.116114504e+00 wpscbe1 = -1.303220350e+02 ppscbe1 = 3.085960190e-5
+ pscbe2 = 2.922546860e-08 lpscbe2 = -9.703471248e-15 wpscbe2 = -6.059420221e-14 ppscbe2 = 2.941550321e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.927406842e+00 lbeta0 = 1.078709509e-08 wbeta0 = 2.723594253e-06 pbeta0 = -8.365991510e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 8.092245841e+08 lbgidl = 1.506150006e+02 wbgidl = 1.630286330e+03 pbgidl = -6.803594825e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.211002050e-01 lkt1 = 1.463071415e-08 wkt1 = 8.318063136e-08 pkt1 = -4.103289036e-14
+ kt2 = -2.863303573e-03 lkt2 = -5.377744449e-09 wkt2 = -1.295510512e-07 pkt2 = 1.310165126e-14
+ at = 1.195361263e+05 lat = -2.202684788e-02 wat = -2.832856651e-01 pat = 7.970835900e-8
+ ute = -4.180238036e-01 lute = 8.358250165e-08 wute = 1.154029435e-06 pute = -2.261081696e-13
+ ua1 = 5.600615966e-09 lua1 = -1.244119505e-15 wua1 = -9.425666971e-15 pua1 = 3.261311382e-21
+ ub1 = -4.469482015e-18 lub1 = 1.057011195e-24 wub1 = 7.846933584e-24 pub1 = -2.892561258e-30
+ uc1 = -7.326917920e-10 luc1 = 1.860693213e-16 wuc1 = 2.154780101e-15 puc1 = -6.337590194e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.286845993e-01 lvth0 = -5.572028975e-08 wvth0 = 6.010354850e-08 pvth0 = 3.887508089e-16
+ k1 = 1.123683124e+00 lk1 = -5.586463061e-08 wk1 = -3.467219483e-06 pk1 = 6.722019082e-13
+ k2 = -1.730916407e-01 lk2 = 1.353098735e-08 wk2 = 1.094355253e-06 pk2 = -2.134662261e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -8.515412636e-01 ldsub = 4.252265561e-07 wdsub = 4.552755307e-06 pdsub = -1.336742769e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.318763268e-01 lvoff = -7.554408177e-09 wvoff = 3.052626130e-07 pvoff = -6.046562781e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -2.541813505e+00 lnfactor = 8.413167520e-07 wnfactor = 1.360503576e-05 pnfactor = -2.255240409e-12
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = -4.195334373e-03 lu0 = 1.896160602e-09 wu0 = 4.922199933e-08 pu0 = -9.819367243e-15
+ ua = -5.413215412e-09 lua = 7.317596187e-16 wua = 1.619518404e-14 pua = -3.167934327e-21
+ ub = 4.702947734e-18 lub = -6.173875712e-25 wub = -1.177555559e-23 pub = 2.352780555e-30
+ uc = 9.989659462e-11 luc = -2.492503702e-17 wuc = -4.460339370e-16 puc = 9.557431995e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.413581281e+04 lvsat = 3.880119724e-03 wvsat = -2.117606890e-01 pvsat = 3.155788742e-8
+ a0 = -3.102288004e-01 la0 = 2.403464363e-07 wa0 = 3.438720520e-06 pa0 = -7.632444697e-13
+ ags = 2.127753980e+00 lags = -1.482263147e-07 wags = 7.847494198e-06 pags = -1.325206345e-12
+ a1 = 0.0
+ a2 = 1.697589778e+00 la2 = -2.144072702e-07 wa2 = -1.726210965e-06 pa2 = 4.123400132e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.356557137e-01 lketa = 9.193296559e-08 wketa = 1.468935435e-06 pketa = -2.901285365e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.980595131e-01 lpclm = -6.248400946e-08 wpclm = -1.496372491e-06 ppclm = 3.589720542e-13
+ pdiblc1 = -8.579017139e-02 lpdiblc1 = 7.685867795e-08 wpdiblc1 = 7.914442929e-07 ppdiblc1 = -8.623582152e-14
+ pdiblc2 = 1.321340355e-02 lpdiblc2 = -9.315706302e-10 wpdiblc2 = -2.951629803e-08 ppdiblc2 = 6.106911695e-15
+ pdiblcb = -2.732510397e-01 lpdiblcb = 5.929972585e-08 wpdiblcb = 2.222728831e-06 ppdiblcb = -5.309432359e-13
+ drout = 1.503710032e+00 ldrout = -2.509636102e-07 wdrout = -5.052048418e-06 pdrout = 1.196103884e-12
+ pscbe1 = 8.029075316e+08 lpscbe1 = -6.409265698e-01 wpscbe1 = -1.038654193e+01 ppscbe1 = 2.210610665e-6
+ pscbe2 = -2.538909488e-08 lpscbe2 = 3.342309529e-15 wpscbe2 = 1.038486722e-13 ppscbe2 = -9.864966207e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.949721164e+00 lbeta0 = 2.443268731e-07 wbeta0 = 6.501395521e-07 pbeta0 = -3.413130265e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.102286019e-10 lagidl = -1.935393061e-16 wagidl = -4.088107259e-15 pagidl = 9.765261809e-22
+ bgidl = 2.166143256e+09 lbgidl = -1.735121626e+02 wbgidl = -3.137448936e+03 pbgidl = 4.585094407e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.962505711e-01 lkt1 = 8.694882115e-09 wkt1 = 2.201926437e-07 pkt1 = -7.376094975e-14
+ kt2 = 5.724519438e-02 lkt2 = -1.973586136e-08 wkt2 = -3.345106921e-07 pkt2 = 6.206036067e-14
+ at = -4.108139137e+04 lat = 1.633985856e-02 wat = 5.085673676e-01 pat = -1.094415749e-7
+ ute = 2.151349326e+00 lute = -5.301636579e-07 wute = -6.405249927e-06 pute = 1.579576892e-12
+ ua1 = 2.175432288e-09 lua1 = -4.259458801e-16 wua1 = 5.606891670e-15 pua1 = -3.295159006e-22
+ ub1 = -2.303763716e-18 lub1 = 5.396860653e-25 wub1 = -4.543604880e-24 pub1 = 6.716666453e-32
+ uc1 = 1.183462596e-10 luc1 = -1.721813812e-17 wuc1 = -1.387329598e-15 puc1 = 2.123447243e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.011847644e+00 lvth0 = -2.728508913e-08 wvth0 = -1.356427282e-07 pvth0 = 3.681124648e-14
+ k1 = -8.773446680e-01 lk1 = 3.104425600e-07 wk1 = 3.635632938e-06 pk1 = -5.803352740e-13
+ k2 = 5.282837761e-01 lk2 = -1.154715083e-07 wk2 = -1.099355141e-06 pk2 = 1.727892604e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.740083934e+00 ldsub = -1.314761622e-06 wdsub = -2.062615595e-05 pdsub = 3.208692702e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.804946298e-02 lvoff = -4.805890324e-08 wvoff = 1.555124573e-07 pvoff = -3.871858994e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.809871638e-01 lnfactor = 2.712284372e-07 wnfactor = -5.308622264e-06 pnfactor = 1.033208064e-12
+ eta0 = 1.893639354e+00 leta0 = -2.608944467e-07 weta0 = -2.169709277e-09 peta0 = 4.032838634e-16
+ etab = 3.394336571e-01 letab = -6.320670259e-08 wetab = -1.038562351e-06 petab = 1.930375841e-13
+ u0 = 2.320625218e-02 lu0 = -3.006087408e-09 wu0 = -4.640976699e-08 pu0 = 6.967201773e-15
+ ua = 3.886184039e-09 lua = -9.230541356e-16 wua = -1.386346346e-14 pua = 2.100153216e-21
+ ub = -2.266581811e-18 lub = 6.158870009e-25 wub = 1.035262472e-23 pub = -1.523331891e-30
+ uc = -2.384631360e-10 luc = 3.545670372e-17 wuc = 7.243663492e-16 puc = -1.123465953e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.330751244e+05 lvsat = -2.713002175e-02 wvsat = -6.722414572e-02 pvsat = 7.869785934e-9
+ a0 = 3.048128637e+00 la0 = -3.596759882e-07 wa0 = -9.225689060e-06 pa0 = 1.513854164e-12
+ ags = 1.25
+ a1 = 0.0
+ a2 = -1.688871825e+00 la2 = 3.934501494e-07 wa2 = 5.608934900e-06 pa2 = -9.095336286e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.688199399e-02 lketa = -1.266460429e-08 wketa = -1.444299522e-06 pketa = 2.221474507e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.075543399e-02 lpclm = 9.243158736e-08 wpclm = 3.822085082e-06 ppclm = -5.934322421e-13
+ pdiblc1 = 1.572835776e+00 lpdiblc1 = -2.236928288e-07 wpdiblc1 = 1.382822590e-06 ppdiblc1 = -2.048365929e-13
+ pdiblc2 = 3.114521763e-02 lpdiblc2 = -4.358337341e-09 wpdiblc2 = 3.613720176e-08 ppdiblc2 = -5.481326679e-15
+ pdiblcb = -5.211727023e+00 lpdiblcb = 9.831839101e-07 wpdiblcb = 2.965908418e-05 ppdiblcb = -5.683988211e-12
+ drout = -5.086777361e+00 ldrout = 9.487459873e-07 wdrout = 1.258301368e-05 pdrout = -1.961314343e-12
+ pscbe1 = 7.944991595e+08 lpscbe1 = 8.574160031e-01 wpscbe1 = 1.675348074e+01 ppscbe1 = -2.611365042e-6
+ pscbe2 = -8.423568013e-08 lpscbe2 = 1.461659180e-14 wpscbe2 = 2.852497637e-13 ppscbe2 = -4.457508489e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.566302834e+01 lbeta0 = -1.164749353e-06 wbeta0 = -6.104997183e-06 pbeta0 = 8.799045449e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.735479305e-09 lagidl = 2.787349843e-16 wagidl = 9.261134760e-15 pagidl = -1.406391369e-21
+ bgidl = 8.467363718e+08 lbgidl = 5.425867241e+01 wbgidl = 4.667830778e+02 pbgidl = -1.652514064e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.940299939e-01 lkt1 = -4.660355016e-08 wkt1 = -6.241926335e-07 pkt1 = 7.575948933e-14
+ kt2 = 3.874109525e-01 lkt2 = -8.309056328e-08 wkt2 = -1.259690573e-06 pkt2 = 2.402711091e-13
+ at = -7.158538946e+04 lat = 2.365455642e-02 wat = 7.076571870e-02 pat = -3.908477318e-8
+ ute = -5.553492691e+00 lute = 8.485642010e-07 wute = 2.095135258e-05 pute = -3.346180148e-12
+ ua1 = -1.307045851e-09 lua1 = 1.784627202e-16 wua1 = 1.346978432e-14 pua1 = -1.824163845e-21
+ ub1 = 9.199194857e-19 lub1 = -5.170191884e-27 wub1 = -9.411370202e-24 pub1 = 9.786998163e-31
+ uc1 = 2.560730738e-11 luc1 = -1.714084476e-18 wuc1 = -1.590789406e-16 puc1 = 5.426338350e-24
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.142549729e+00 lvth0 = 1.077794445e-06 wvth0 = 8.424617286e-08 pvth0 = -1.683985797e-12
+ k1 = 4.303698969e-01 lk1 = 1.109590230e-06 wk1 = -1.863414147e-08 pk1 = 3.724754314e-13
+ k2 = 2.209900758e-02 lk2 = -2.409044937e-07 wk2 = 3.082242674e-08 pk2 = -6.161054813e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.787253552e-01 lvoff = -1.281417789e-06 wvoff = -1.186857965e-07 pvoff = 2.372394957e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 4.130185353e+00 lnfactor = -5.166596095e-05 wnfactor = -5.191106049e-06 pnfactor = 1.037643440e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.510124600e-02 lu0 = -4.409891208e-07 wu0 = -4.218960189e-08 pu0 = 8.433224676e-13
+ ua = 7.053534227e-10 lua = -2.629029356e-14 wua = -2.736587223e-15 pua = 5.470128624e-20
+ ub = 3.831042496e-18 lub = -4.327535737e-23 wub = -4.013641232e-24 pub = 8.022815281e-29
+ uc = -6.496972548e-11 luc = -8.841609808e-16 wuc = -1.468731067e-17 puc = 2.935827436e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.113870874e+05 lvsat = -3.019810289e+00 wvsat = -3.090414997e-01 pvsat = 6.177390362e-6
+ a0 = 1.165770398e+00 la0 = 9.067415208e-06 wa0 = 9.337106358e-07 pa0 = -1.866382052e-11
+ ags = 1.039916176e-01 lags = 7.515813769e-06 wags = 7.738276898e-07 pags = -1.546794109e-11
+ a1 = 0.0
+ a2 = 1.561282690e+00 la2 = -1.521718071e-05 wa2 = -1.557296618e-06 pa2 = 3.112859965e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = 8.574671297e-02 lketa = -2.338351742e-06 wketa = -2.875115450e-07 pketa = 5.747030896e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.762746415e-01 lpclm = 4.725784767e-06 wpclm = 7.784550232e-07 ppclm = -1.556043626e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.331171642e-02 lpdiblc2 = -2.603495722e-07 wpdiblc2 = -2.695201662e-08 ppdiblc2 = 5.387403565e-13
+ pdiblcb = 7.855039219e-03 lpdiblcb = -1.876027773e-07 wpdiblcb = -2.312339226e-08 ppdiblcb = 4.622104819e-13
+ drout = 0.56
+ pscbe1 = 8.064388516e+08 lpscbe1 = -3.234049569e+02 wpscbe1 = -2.159460135e+02 ppscbe1 = 4.316516791e-3
+ pscbe2 = 9.285602072e-09 lpscbe2 = 1.497834542e-15 wpscbe2 = 7.781094574e-16 ppscbe2 = -1.555352879e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.576215346e-10 lalpha0 = 1.914177236e-14 walpha0 = 2.916553213e-15 palpha0 = -5.829860303e-20
+ alpha1 = 3.549704974e-10 lalpha1 = -5.096572126e-15 walpha1 = -7.765437562e-16 palpha1 = 1.552223219e-20
+ beta0 = 9.273771998e+00 lbeta0 = -1.254056129e-04 wbeta0 = -1.228462290e-05 pbeta0 = 2.455557302e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.852343277e-11 lagidl = 1.147528989e-15
+ bgidl = 4.363286167e+08 lbgidl = 1.126715400e+04 wbgidl = 2.304639364e+03 pbgidl = -4.606713664e-2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.637968559e-01 lkt1 = 1.650452194e-07 wkt1 = 7.786872433e-08 pkt1 = -1.556507808e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -1.653904217e-01 lute = -3.284162913e-06 wute = -3.898887027e-07 pute = 7.793434593e-12
+ ua1 = 2.139764998e-09 lua1 = 7.182700633e-15
+ ub1 = -2.472812867e-19 lub1 = -2.865441920e-23 wub1 = -9.886991928e-25 pub1 = 1.976297963e-29
+ uc1 = 4.338507642e-11 luc1 = 7.645641303e-15 puc1 = -3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.08863
+ k1 = 0.4858803
+ k2 = 0.010047076
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.24283192
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.5454489
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0130395126
+ ua = -6.0989319e-10
+ ub = 1.66606982e-18
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.6193936
+ ags = 0.47999155
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.093872372e+00 lvth0 = 4.188063158e-8
+ k1 = 4.522972755e-01 lk1 = 2.682904169e-7
+ k2 = 2.243897693e-02 lk2 = -9.899728555e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.402497948e-01 lvoff = -2.062826246e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.707115507e+00 lnfactor = -1.291533511e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.609958679e-02 lu0 = -2.444653486e-8
+ ua = -1.211989359e-10 lua = -3.904114865e-15
+ ub = 1.642518584e-18 lub = 1.881477614e-25
+ uc = -1.423307551e-10 luc = 2.646582022e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.212579461e+05 lvsat = -4.868852462e-1
+ a0 = 1.674871402e+00 la0 = -4.432049504e-7
+ ags = 4.562623108e-01 lags = 1.895698069e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.743565127e-02 lketa = 4.952840774e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.109267259e-01 lpclm = 4.562227086e-06 wpclm = 1.110223025e-22 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.587787891e-04 lpdiblc2 = -5.735148984e-10
+ pdiblcb = -4.459427061e-04 lpdiblcb = -8.662970003e-9
+ drout = 0.56
+ pscbe1 = 7.805463027e+08 lpscbe1 = 7.759826970e+1
+ pscbe2 = 9.153007757e-09 lpscbe2 = 1.657912159e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.819567689e-01 lbeta0 = 2.941467397e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.917358547e-10 lagidl = -3.659223987e-16
+ bgidl = 8.022575536e+08 lbgidl = 1.579738698e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.101376581e-01 lkt1 = 4.361735931e-7
+ kt2 = -3.138933667e-02 lkt2 = -5.250016399e-8
+ at = -1.789107917e+05 lat = 1.429295056e+0
+ ute = 1.617288118e-01 lute = -3.925881003e-6
+ ua1 = 5.328096354e-09 lua1 = -2.260048410e-14
+ ub1 = -4.224512371e-18 lub1 = 2.032138745e-23
+ uc1 = 7.901037197e-10 luc1 = -2.909735948e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.091123626e+00 lvth0 = 3.091624109e-8
+ k1 = 5.977558582e-01 lk1 = -3.119249599e-7
+ k2 = -2.975396524e-02 lk2 = 1.091935757e-07 wk2 = 3.469446952e-24 pk2 = -6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.223229514e-01 lvoff = -9.213611045e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.717805832e+00 lnfactor = -1.334175826e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.150387845e-03 lu0 = 7.261786318e-9
+ ua = -1.665485757e-09 lua = 2.255844507e-15
+ ub = 2.098150966e-18 lub = -1.629310578e-24
+ uc = -6.694967090e-11 luc = -3.602714318e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.447013512e+05 lvsat = -1.815109412e-1
+ a0 = 1.964115559e+00 la0 = -1.596962289e-6
+ ags = 6.423764338e-01 lags = -5.528152347e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.118284482e-02 lketa = 6.447547569e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.336218480e-01 lpclm = -1.199889384e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 1.963998626e-02 lpdiblcb = -8.878312947e-08 wpdiblcb = -6.938893904e-24 ppdiblcb = 1.387778781e-29
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.671893803e-08 lpscbe2 = -2.852160011e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.565947440e+00 lbeta0 = 4.492596311e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.143013757e+09 lbgidl = 2.205064997e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.434839429e-01 lkt1 = -2.285864121e-7
+ kt2 = -4.017360155e-02 lkt2 = -1.746087337e-8
+ at = 2.745973838e+05 lat = -3.796900997e-1
+ ute = -1.640382899e+00 lute = 3.262508336e-6
+ ua1 = -3.274541222e-09 lua1 = 1.171431885e-14 wua1 = -8.271806126e-31 pua1 = -1.654361225e-36
+ ub1 = 3.170152177e-18 lub1 = -9.174968124e-24
+ uc1 = 9.216446460e-11 luc1 = -1.257469911e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.090838253e+00 lvth0 = 3.034867045e-8
+ k1 = 4.322967437e-01 lk1 = 1.715170913e-8
+ k2 = 2.844424485e-02 lk2 = -6.555098444e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.916658762e-01 ldsub = 3.347946888e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.996927125e-01 lvoff = 6.174228629e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.177495674e-01 lnfactor = 1.649241077e-6
+ eta0 = -5.744849986e-02 leta0 = 2.733671979e-07 peta0 = 1.110223025e-28
+ etab = 6.842919891e-01 letab = -1.500188708e-06 wetab = -3.330669074e-22 petab = -1.110223025e-28
+ u0 = 1.359283912e-02 lu0 = -3.562541745e-9
+ ua = -1.917591780e-10 lua = -6.752060745e-16
+ ub = 1.151418582e-18 lub = 2.536170597e-25
+ uc = -1.214437714e-10 luc = 7.235453841e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.038194939e+04 lvsat = 2.596678738e-2
+ a0 = 1.115812466e+00 la0 = 9.020228253e-8
+ ags = 1.549979248e-01 lags = 4.165172605e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.629453859e-03 lketa = -1.220220699e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.108255342e-02 lpclm = 5.752552428e-7
+ pdiblc1 = 4.088045794e-01 lpdiblc1 = -3.739986375e-8
+ pdiblc2 = 2.392950000e-06 lpdiblc2 = 4.228477835e-10
+ pdiblcb = -0.025
+ drout = 1.344068365e-01 ldrout = 8.464494752e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.454152232e-09 lpscbe2 = 1.358892391e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.794355910e+00 lbeta0 = 2.049451557e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.269088568e+09 lbgidl = -3.023991007e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444605805e-01 lkt1 = -2.775700689e-8
+ kt2 = -6.040588351e-02 lkt2 = 2.277850526e-8
+ at = 6.493100483e+04 lat = 3.730907145e-2
+ ute = 0.0
+ ua1 = 2.824339679e-09 lua1 = -4.155624112e-16
+ ub1 = -1.527062104e-18 lub1 = 1.671804431e-25
+ uc1 = 1.528486051e-10 luc1 = -2.464398577e-16 wuc1 = -5.169878828e-32 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.083811263e+00 lvth0 = 2.339989136e-8
+ k1 = 3.328536151e-01 lk1 = 1.154880357e-7
+ k2 = 6.118412774e-02 lk2 = -3.893058644e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.664626476e-01 ldsub = 2.608304055e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.329295969e-01 lvoff = -4.277755777e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.557974615e+00 lnfactor = 3.239327345e-7
+ eta0 = 3.582529886e-01 leta0 = -1.377075330e-7
+ etab = -1.646537114e+00 letab = 8.046982669e-7
+ u0 = 1.168706777e-02 lu0 = -1.677981632e-9
+ ua = -5.906662208e-10 lua = -2.807388671e-16
+ ub = 1.291920204e-18 lub = 1.146792206e-25
+ uc = -6.422249855e-11 luc = 1.577013837e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.500133002e+04 lvsat = 1.621420453e-3
+ a0 = 1.232969442e+00 la0 = -2.565073621e-8
+ ags = -8.543032923e-02 lags = 6.542695481e-07 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 6.044617774e-01 la2 = 1.933618822e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.631183582e-02 lketa = -3.093268012e-08 pketa = -1.387778781e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.378830106e-01 lpclm = 8.398417474e-8
+ pdiblc1 = -2.440305587e-01 lpdiblc1 = 6.081692192e-7
+ pdiblc2 = -1.444786656e-04 lpdiblc2 = 5.680847180e-10
+ pdiblcb = -4.911716338e-02 lpdiblcb = 2.384873935e-8
+ drout = 1.009114736e+00 ldrout = -1.852292549e-8
+ pscbe1 = 8.085510012e+08 lpscbe1 = -8.455828520e+0
+ pscbe2 = 9.336779542e-09 lpscbe2 = -4.851479500e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.461134792e+00 lbeta0 = 4.012239235e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.280411890e+09 lbgidl = -4.143720287e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.540604914e-01 lkt1 = -1.826394297e-8
+ kt2 = -2.736871980e-02 lkt2 = -9.890954821e-9
+ at = 1.688138884e+05 lat = -6.541759562e-2
+ ute = 1.955480000e-02 lute = -1.933715508e-8
+ ua1 = 2.651272672e-09 lua1 = -2.444216402e-16 wua1 = -3.308722450e-30
+ ub1 = -1.049425256e-18 lub1 = -3.051403071e-25
+ uc1 = -1.219162794e-10 luc1 = 2.526689368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.030465367e+00 lvth0 = -2.679317192e-9
+ k1 = 4.675435820e-01 lk1 = 4.964215164e-8
+ k2 = 1.221796632e-02 lk2 = -1.499249910e-08 pk2 = 6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.395528179e+00 ldsub = -1.933618609e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.371839266e-01 lvoff = -2.197941611e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.099442871e+00 lnfactor = 5.922514810e-8
+ eta0 = -3.184587778e-01 leta0 = 1.931165483e-07 peta0 = 5.551115123e-29
+ etab = -3.801533128e-04 letab = -5.848652817e-11
+ u0 = 1.002014040e-02 lu0 = -8.630708464e-10
+ ua = -9.529635079e-10 lua = -1.036225924e-16
+ ub = 1.565225622e-18 lub = -1.893159938e-26
+ uc = -4.384699617e-11 luc = 5.809166520e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.178071320e+04 lvsat = -6.581516602e-3
+ a0 = 1.567087208e+00 la0 = -1.889908884e-7
+ ags = 2.884384880e-01 lags = 4.714962994e-7
+ a1 = 0.0
+ a2 = 1.191076445e+00 la2 = -9.341643046e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.755142380e-02 lketa = -9.489248387e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.776001892e-01 lpclm = -3.320636238e-8
+ pdiblc1 = 1.594980969e+00 lpdiblc1 = -2.908683466e-7
+ pdiblc2 = -5.669698530e-03 lpdiblc2 = 3.269198953e-9
+ pdiblcb = 2.323432675e-02 lpdiblcb = -1.152173363e-08 wpdiblcb = -9.540979118e-24 ppdiblcb = -6.396792818e-30
+ drout = 1.480326837e+00 ldrout = -2.488843850e-7
+ pscbe1 = 7.830387781e+08 lpscbe1 = 4.016331970e+0
+ pscbe2 = 9.329958843e-09 lpscbe2 = -4.518035983e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.821672202e+00 lbeta0 = -2.639019999e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.344513051e+09 lbgidl = -7.277433743e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.937886636e-01 lkt1 = 1.157968567e-9
+ kt2 = -4.540011584e-02 lkt2 = -1.075946241e-9
+ at = 2.652206705e+04 lat = 4.144607083e-3
+ ute = -3.910960000e-02 lute = 9.342110152e-9
+ ua1 = 2.505791010e-09 lua1 = -1.733000203e-16
+ ub1 = -1.893018625e-18 lub1 = 1.072671831e-25
+ uc1 = -2.519095944e-11 luc1 = -2.201921350e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.089501693e-01 lvth0 = -5.559265240e-08 wvth0 = -6.569671029e-14 pvth0 = 1.569297314e-20
+ k1 = -1.474413380e-02 lk1 = 1.648462183e-07 wk1 = -3.816552709e-13 pk1 = 9.116599431e-20
+ k2 = 1.862291287e-01 lk2 = -5.655854547e-08 wk2 = 1.250127735e-14 pk2 = -2.986180192e-21
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.433110956e-01 ldsub = -1.367976616e-08 wdsub = 7.455866324e-14 pdsub = -1.780982783e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.316463403e-01 lvoff = -2.740770487e-08 wvoff = -3.922896408e-14 pvoff = 9.370622722e-21
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.925266402e+00 lnfactor = 1.008306812e-07 wnfactor = -1.085649657e-12 pnfactor = 2.593291342e-19
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 1.196622625e-02 lu0 = -1.327932374e-09 wu0 = -5.246282880e-15 pu0 = 1.253179595e-21
+ ua = -9.568609602e-11 lua = -3.084004478e-16 wua = -2.315927408e-22 pua = 5.532055806e-29
+ ub = 8.365600827e-19 lub = 1.551247380e-25 wub = -2.955879191e-31 pub = 7.060708546e-38
+ uc = -4.655425743e-11 luc = 6.455850017e-18 wuc = -7.089599594e-26 puc = 1.693493330e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.393735735e+03 lvsat = 1.424184401e-02 wvsat = 3.365099546e-08 pvsat = -8.038213244e-15
+ a0 = 8.188412249e-01 la0 = -1.025737040e-08 wa0 = 1.110700154e-14 pa0 = -2.653129272e-21
+ ags = 4.704401308e+00 lags = -5.833447395e-07 wags = 4.100134916e-13 pags = -9.793992106e-20
+ a1 = 0.0
+ a2 = 1.130805108e+00 la2 = -7.901941609e-08 wa2 = 8.951765587e-13 pa2 = -2.138308242e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.334522481e-02 lketa = -3.327883141e-09 wketa = -5.907980771e-16 pketa = 1.411240014e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.067403384e-01 lpclm = 5.538093019e-08 wpclm = -3.899264911e-15 ppclm = 9.314176097e-22
+ pdiblc1 = 1.740727862e-01 lpdiblc1 = 4.854399118e-08 wpdiblc1 = -4.785460561e-14 ppdiblc1 = 1.143102946e-20
+ pdiblc2 = 3.522017863e-03 lpdiblc2 = 1.073573658e-09 wpdiblc2 = -5.742553377e-16 ppdiblc2 = 1.371723707e-22
+ pdiblcb = 4.565600017e-01 lpdiblcb = -1.150302376e-07 wpdiblcb = 2.677494785e-13 ppdiblcb = -6.395731800e-20
+ drout = -1.550803608e-01 ldrout = 1.417653322e-07 wdrout = 9.618185182e-14 pdrout = -2.297495882e-20
+ pscbe1 = 7.994972153e+08 lpscbe1 = 8.490506716e-02 wpscbe1 = -7.798528671e-06 ppscbe1 = 1.862834930e-12
+ pscbe2 = 8.708594014e-09 lpscbe2 = 1.032450570e-16 wpscbe2 = 7.999399536e-22 ppscbe2 = -1.910816596e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.163187944e+00 lbeta0 = 1.322601349e-07 wbeta0 = 4.312823023e-13 pbeta0 = -1.030204047e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.320611150e-10 lagidl = 1.270934385e-16 wagidl = -1.666049370e-22 pagidl = 3.979692119e-29
+ bgidl = 1.135992664e+09 lbgidl = -2.296507275e+01 wbgidl = 3.698393135e-04 pbgidl = -8.834351635e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.239524495e-01 lkt1 = -1.552380789e-08 wkt1 = -1.061072474e-13 pkt1 = 2.534583832e-20
+ kt2 = -5.258809566e-02 lkt2 = 6.410464987e-10 wkt2 = -7.603565111e-15 pkt2 = 1.816263584e-21
+ at = 1.259016779e+05 lat = -1.959420056e-02 wat = 5.825264635e-08 pat = -1.391480965e-14
+ ute = 4.824857555e-02 lute = -1.152513724e-08 wute = -1.254854221e-14 pute = 2.997470272e-21
+ ua1 = 4.016400244e-09 lua1 = -5.341392479e-16 wua1 = -8.401142233e-22 pua1 = 2.006780839e-28
+ ub1 = -3.795611892e-18 lub1 = 5.617396367e-25 wub1 = 7.444050248e-31 pub1 = -1.778160289e-37
+ uc1 = -3.371697339e-10 luc1 = 5.250315636e-17 wuc1 = -6.676013217e-23 puc1 = 1.594699272e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.056384299e+00 lvth0 = -1.519853600e-08 wvth0 = -9.108421537e-13 pvth0 = 1.743599531e-19
+ k1 = 3.163794938e-01 lk1 = 1.198951989e-07 wk1 = 3.685256118e-13 pk1 = -3.909252211e-20
+ k2 = 1.673213808e-01 lk2 = -5.873786326e-08 wk2 = -1.282034932e-13 pk2 = 2.286599943e-20
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.967688838e+00 ldsub = -2.612189876e-07 wdsub = -4.483775840e-13 pdsub = 7.759543186e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.301151156e-02 lvoff = -6.077177024e-08 wvoff = 2.986523207e-14 pvoff = -2.528582899e-21
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -7.620475502e-01 lnfactor = 6.104722649e-07 wnfactor = 2.607350538e-12 pnfactor = -4.009823691e-19
+ eta0 = 1.892926871e+00 leta0 = -2.607620175e-07 weta0 = 2.447968441e-13 peta0 = -4.550038968e-20
+ etab = -1.568066564e-03 letab = 1.752877822e-10 wetab = 8.391869422e-16 petab = -1.559796775e-22
+ u0 = 7.968055921e-03 lu0 = -7.184742834e-10 wu0 = 1.877871497e-14 pu0 = -3.086190224e-21
+ ua = -6.657480479e-10 lua = -2.334894449e-16 wua = 1.045366863e-21 pua = -1.764588485e-28
+ ub = 1.132600365e-18 lub = 1.157160070e-25 wub = 7.047681971e-31 pub = -1.082211513e-37
+ uc = -6.245784946e-13 luc = -1.431194449e-18 wuc = 6.015200804e-24 puc = -1.112583075e-30
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.110028048e+05 lvsat = -2.454606659e-02 wvsat = -2.037378815e-07 pvsat = 3.527605708e-14
+ a0 = 1.896421654e-02 la0 = 1.373831684e-07 wa0 = 7.414769492e-13 pa0 = -1.386740793e-19
+ ags = 1.250000346e+00 lags = -5.389125057e-14 wags = -1.053008134e-12 pags = 1.641323779e-19
+ a1 = 0.0
+ a2 = 1.527674086e-01 la2 = 9.481363330e-08 wa2 = -2.065570250e-12 pa2 = 3.149570160e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.973396729e-01 lketa = 6.027534974e-08 wketa = 4.199554233e-13 pketa = -7.801159535e-20
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.285699180e+00 lpclm = -1.024159983e-07 wpclm = 8.004728080e-13 ppclm = -1.484834549e-19
+ pdiblc1 = 2.026872356e+00 lpdiblc1 = -2.909489823e-07 wpdiblc1 = -1.206082928e-12 ppdiblc1 = 2.278616802e-19
+ pdiblc2 = 4.301049316e-02 lpdiblc2 = -6.158073494e-09 wpdiblc2 = 5.757148719e-14 ppdiblc2 = -1.065656776e-20
+ pdiblcb = 4.526545287e+00 lpdiblcb = -8.830983993e-07 wpdiblcb = -1.221049108e-11 ppdiblcb = 2.248934727e-18
+ drout = -9.552692295e-01 ldrout = 3.047678332e-07 wdrout = 1.623279807e-12 pdrout = -3.091295264e-19
+ pscbe1 = 7.999999934e+08 lpscbe1 = 1.025021076e-06 wpscbe1 = 2.002840424e-05 ppscbe1 = -3.121827126e-12
+ pscbe2 = 9.423272207e-09 lpscbe2 = -1.919858632e-17 wpscbe2 = -1.991224164e-21 ppscbe2 = 3.084759924e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.365851252e+01 lbeta0 = -8.758413281e-07 wbeta0 = 3.080038482e-13 pbeta0 = -9.047761296e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.305323381e-09 lagidl = -1.830398288e-16 wagidl = -7.961726653e-22 pagidl = 1.608209977e-28
+ bgidl = 1.000000312e+09 lbgidl = -4.861084700e-05 wbgidl = -9.498316803e-04 pbgidl = 1.480502644e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.989776034e-01 lkt1 = -2.172865114e-08 wkt1 = 3.149834562e-13 pkt1 = -5.037074624e-20
+ kt2 = -2.619607966e-02 lkt2 = -4.199903906e-09 wkt2 = 1.035279331e-13 pkt2 = -1.865690624e-20
+ at = -4.835015559e+04 lat = 1.082145614e-02 wat = -2.075133112e-08 pat = -6.311324396e-16
+ ute = 1.325677818e+00 lute = -2.501211363e-07 wute = -4.604924002e-13 pute = 8.655854808e-20
+ ua1 = 3.115624181e-09 lua1 = -4.204833471e-16 wua1 = 3.175666108e-21 pua1 = -5.255329125e-28
+ ub1 = -2.170210357e-18 lub1 = 3.161761073e-25 wub1 = -2.771513092e-30 pub1 = 4.577870828e-37
+ uc1 = -2.662475279e-11 luc1 = 6.760904313e-20 wuc1 = 1.709455309e-22 puc1 = -2.662998859e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.101366082e+00 lvth0 = 2.545798937e-7
+ k1 = 4.212606180e-01 lk1 = 1.291674424e-6
+ k2 = 3.716651602e-02 lk2 = -5.420869610e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.367447726e-01 lvoff = -1.216751986e-07 wvoff = 4.440892099e-22
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.592519036e+00 lnfactor = -9.408788196e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.447690685e-02 lu0 = -2.873188681e-8
+ ua = -6.324241445e-10 lua = 4.503683210e-16
+ ub = 1.868978521e-18 lub = -4.055915651e-24 wub = -3.081487911e-39
+ uc = -7.214960068e-11 luc = -7.406433888e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.622213786e+00 la0 = -5.637233290e-8
+ ags = 4.822764082e-01 lags = -4.567173287e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.480298045e-02 lketa = 4.710778082e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.042722157e-01 lpclm = -2.880916892e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.362535913e-04 lpdiblc2 = 3.013041483e-9
+ pdiblcb = -3.448804924e-03 lpdiblcb = 3.834829377e-8
+ drout = 0.56
+ pscbe1 = 7.008738872e+08 lpscbe1 = 1.786719392e+3
+ pscbe2 = 9.665980000e-09 lpscbe2 = -6.105490408e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.681322036e-10 lalpha0 = -9.357433760e-15
+ alpha1 = -2.464203913e-11 lalpha1 = 2.491453517e-15 palpha1 = -2.197198502e-37
+ beta0 = 3.268447993e+00 lbeta0 = -5.365972042e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.852343277e-11 lagidl = 1.147528989e-15
+ bgidl = 1.562948962e+09 lbgidl = -1.125271361e+4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.257308181e-01 lkt1 = -5.958518612e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.559870728e-01 lute = 5.256487698e-7
+ ua1 = 2.139764998e-09 lua1 = 7.182700633e-15
+ ub1 = -7.306057684e-19 lub1 = -1.899330897e-23
+ uc1 = 4.338507642e-11 luc1 = 7.645641303e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.08863
+ k1 = 0.4858803
+ k2 = 0.010047076
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.24283192
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.5454489
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0130395126
+ ua = -6.0989319e-10
+ ub = 1.66606982e-18
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.6193936
+ ags = 0.47999155
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.093872372e+00 lvth0 = 4.188063158e-8
+ k1 = 4.522972755e-01 lk1 = 2.682904169e-7
+ k2 = 2.243897693e-02 lk2 = -9.899728555e-08 pk2 = 1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.402497948e-01 lvoff = -2.062826246e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.707115507e+00 lnfactor = -1.291533511e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.609958679e-02 lu0 = -2.444653486e-8
+ ua = -1.211989359e-10 lua = -3.904114865e-15
+ ub = 1.642518584e-18 lub = 1.881477614e-25
+ uc = -1.423307551e-10 luc = 2.646582022e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.212579461e+05 lvsat = -4.868852462e-1
+ a0 = 1.674871402e+00 la0 = -4.432049504e-7
+ ags = 4.562623108e-01 lags = 1.895698069e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.743565127e-02 lketa = 4.952840774e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.109267259e-01 lpclm = 4.562227086e-06 wpclm = -4.440892099e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 3.587787891e-04 lpdiblc2 = -5.735148984e-10
+ pdiblcb = -4.459427061e-04 lpdiblcb = -8.662970003e-9
+ drout = 0.56
+ pscbe1 = 7.805463027e+08 lpscbe1 = 7.759826970e+1
+ pscbe2 = 9.153007757e-09 lpscbe2 = 1.657912159e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.819567689e-01 lbeta0 = 2.941467397e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.917358547e-10 lagidl = -3.659223987e-16
+ bgidl = 8.022575536e+08 lbgidl = 1.579738698e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.101376581e-01 lkt1 = 4.361735931e-7
+ kt2 = -3.138933667e-02 lkt2 = -5.250016399e-8
+ at = -1.789107917e+05 lat = 1.429295056e+0
+ ute = 1.617288118e-01 lute = -3.925881003e-6
+ ua1 = 5.328096354e-09 lua1 = -2.260048410e-14 pua1 = -2.646977960e-35
+ ub1 = -4.224512371e-18 lub1 = 2.032138745e-23 pub1 = 2.465190329e-44
+ uc1 = 7.901037197e-10 luc1 = -2.909735948e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.091123626e+00 lvth0 = 3.091624109e-8
+ k1 = 5.977558582e-01 lk1 = -3.119249599e-7
+ k2 = -2.975396524e-02 lk2 = 1.091935757e-07 wk2 = 2.081668171e-23 pk2 = -1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.223229514e-01 lvoff = -9.213611045e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.717805832e+00 lnfactor = -1.334175826e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.150387845e-03 lu0 = 7.261786318e-9
+ ua = -1.665485757e-09 lua = 2.255844507e-15
+ ub = 2.098150966e-18 lub = -1.629310578e-24
+ uc = -6.694967090e-11 luc = -3.602714318e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.447013512e+05 lvsat = -1.815109412e-1
+ a0 = 1.964115559e+00 la0 = -1.596962289e-6
+ ags = 6.423764338e-01 lags = -5.528152347e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.118284482e-02 lketa = 6.447547569e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.336218480e-01 lpclm = -1.199889384e-06 wpclm = 1.776356839e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 1.963998626e-02 lpdiblcb = -8.878312947e-08 ppdiblcb = -4.163336342e-29
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.671893803e-08 lpscbe2 = -2.852160011e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.565947440e+00 lbeta0 = 4.492596311e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.143013757e+09 lbgidl = 2.205064997e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.434839429e-01 lkt1 = -2.285864121e-7
+ kt2 = -4.017360155e-02 lkt2 = -1.746087337e-8
+ at = 2.745973838e+05 lat = -3.796900997e-1
+ ute = -1.640382899e+00 lute = 3.262508336e-6
+ ua1 = -3.274541222e-09 lua1 = 1.171431885e-14 wua1 = 8.271806126e-31 pua1 = 8.271806126e-36
+ ub1 = 3.170152177e-18 lub1 = -9.174968124e-24 wub1 = 3.081487911e-39 pub1 = 6.162975822e-45
+ uc1 = 9.216446460e-11 luc1 = -1.257469911e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.090838253e+00 lvth0 = 3.034867045e-8
+ k1 = 4.322967437e-01 lk1 = 1.715170913e-8
+ k2 = 2.844424485e-02 lk2 = -6.555098444e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.916658762e-01 ldsub = 3.347946888e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.996927125e-01 lvoff = 6.174228629e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.177495674e-01 lnfactor = 1.649241077e-6
+ eta0 = -5.744849986e-02 leta0 = 2.733671979e-7
+ etab = 6.842919891e-01 letab = -1.500188708e-06 wetab = 2.220446049e-22 petab = -1.554312234e-27
+ u0 = 1.359283912e-02 lu0 = -3.562541745e-9
+ ua = -1.917591780e-10 lua = -6.752060745e-16
+ ub = 1.151418582e-18 lub = 2.536170597e-25
+ uc = -1.214437714e-10 luc = 7.235453841e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.038194939e+04 lvsat = 2.596678738e-2
+ a0 = 1.115812466e+00 la0 = 9.020228253e-8
+ ags = 1.549979248e-01 lags = 4.165172605e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.629453859e-03 lketa = -1.220220699e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.108255342e-02 lpclm = 5.752552428e-7
+ pdiblc1 = 4.088045794e-01 lpdiblc1 = -3.739986375e-8
+ pdiblc2 = 2.392950000e-06 lpdiblc2 = 4.228477835e-10
+ pdiblcb = -0.025
+ drout = 1.344068365e-01 ldrout = 8.464494752e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.454152232e-09 lpscbe2 = 1.358892391e-14 ppscbe2 = 1.323488980e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.794355910e+00 lbeta0 = 2.049451557e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.269088568e+09 lbgidl = -3.023991007e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444605805e-01 lkt1 = -2.775700689e-8
+ kt2 = -6.040588351e-02 lkt2 = 2.277850526e-8
+ at = 6.493100483e+04 lat = 3.730907145e-2
+ ute = 0.0
+ ua1 = 2.824339679e-09 lua1 = -4.155624112e-16
+ ub1 = -1.527062104e-18 lub1 = 1.671804431e-25
+ uc1 = 1.528486051e-10 luc1 = -2.464398577e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.083811263e+00 lvth0 = 2.339989136e-8
+ k1 = 3.328536151e-01 lk1 = 1.154880357e-7
+ k2 = 6.118412774e-02 lk2 = -3.893058644e-08 pk2 = 2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.664626476e-01 ldsub = 2.608304055e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.329295969e-01 lvoff = -4.277755777e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.557974615e+00 lnfactor = 3.239327345e-7
+ eta0 = 3.582529886e-01 leta0 = -1.377075330e-7
+ etab = -1.646537114e+00 letab = 8.046982669e-7
+ u0 = 1.168706777e-02 lu0 = -1.677981632e-9
+ ua = -5.906662208e-10 lua = -2.807388671e-16
+ ub = 1.291920204e-18 lub = 1.146792206e-25
+ uc = -6.422249855e-11 luc = 1.577013837e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.500133002e+04 lvsat = 1.621420453e-3
+ a0 = 1.232969442e+00 la0 = -2.565073621e-8
+ ags = -8.543032923e-02 lags = 6.542695481e-7
+ a1 = 0.0
+ a2 = 6.044617774e-01 la2 = 1.933618822e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.631183582e-02 lketa = -3.093268012e-08 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.378830106e-01 lpclm = 8.398417474e-8
+ pdiblc1 = -2.440305587e-01 lpdiblc1 = 6.081692192e-7
+ pdiblc2 = -1.444786656e-04 lpdiblc2 = 5.680847180e-10
+ pdiblcb = -4.911716338e-02 lpdiblcb = 2.384873935e-8
+ drout = 1.009114736e+00 ldrout = -1.852292549e-8
+ pscbe1 = 8.085510012e+08 lpscbe1 = -8.455828520e+0
+ pscbe2 = 9.336779542e-09 lpscbe2 = -4.851479500e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.461134792e+00 lbeta0 = 4.012239235e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.280411890e+09 lbgidl = -4.143720287e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.540604914e-01 lkt1 = -1.826394297e-8
+ kt2 = -2.736871980e-02 lkt2 = -9.890954821e-9
+ at = 1.688138884e+05 lat = -6.541759562e-2
+ ute = 1.955480000e-02 lute = -1.933715508e-8
+ ua1 = 2.651272672e-09 lua1 = -2.444216402e-16
+ ub1 = -1.049425256e-18 lub1 = -3.051403071e-25
+ uc1 = -1.219162794e-10 luc1 = 2.526689368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.527536513e+00 lvth0 = 2.403238540e-07 wvth0 = 1.016819672e-06 pvth0 = -4.970926330e-13
+ k1 = 1.941485345e+00 lk1 = -6.709237583e-07 wk1 = -3.015127698e-06 pk1 = 1.474005478e-12
+ k2 = -4.934896120e-01 lk2 = 2.322327647e-07 wk2 = 1.034486548e-06 pk2 = -5.057294386e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.273213053e+00 ldsub = -1.335656650e-07 wdsub = 2.502105136e-07 pdsub = -1.223204138e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -4.822447087e-01 lvoff = 1.176049229e-07 wvoff = 5.013017271e-07 pvoff = -2.450713753e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.001002520e+00 lnfactor = -3.815203175e-07 wnfactor = -1.844250252e-06 pnfactor = 9.015986208e-13
+ eta0 = -3.184587778e-01 leta0 = 1.931165483e-07 weta0 = 2.220446049e-22 peta0 = 2.220446049e-28
+ etab = -3.801533128e-04 letab = -5.848652817e-11
+ u0 = -1.853310949e-03 lu0 = 4.941503312e-09 wu0 = 2.428859329e-08 pu0 = -1.187396460e-14
+ ua = -3.710467694e-09 lua = 1.244438479e-15 wua = 5.640811229e-15 pua = -2.757623385e-21
+ ub = 2.952244514e-18 lub = -6.970035250e-25 wub = -2.837316359e-24 pub = 1.387078849e-30
+ uc = 1.387676902e-11 luc = -2.241025057e-17 wuc = -1.180810040e-16 puc = 5.772626043e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.091214398e+05 lvsat = -6.883457761e-02 wvsat = -2.604909918e-01 pvsat = 1.273462312e-7
+ a0 = 1.475372854e+00 la0 = -1.441544921e-07 wa0 = 1.876129005e-07 pa0 = -9.171831865e-14
+ ags = -4.927428888e+00 lags = 3.021377384e-06 wags = 1.066969305e-05 pags = -5.216092843e-12
+ a1 = 0.0
+ a2 = 4.845383075e-01 la2 = 2.519888689e-07 wa2 = 1.445309958e-06 pa2 = -7.065686794e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.730706253e-02 lketa = 5.057390717e-09 wketa = 6.086878920e-08 pketa = -2.975692498e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.272778334e+00 lpclm = -2.752841019e-07 wpclm = -1.012947306e-06 ppclm = 4.951995497e-13
+ pdiblc1 = 2.029027959e+00 lpdiblc1 = -5.030608985e-07 wpdiblc1 = -8.878960716e-07 ppdiblc1 = 4.340657525e-13
+ pdiblc2 = 3.929458420e-03 lpdiblc2 = -1.423540905e-09 wpdiblc2 = -1.963624664e-08 ppdiblc2 = 9.599571893e-15
+ pdiblcb = -1.005287123e+00 lpdiblcb = 4.912915477e-07 wpdiblcb = 2.103966106e-06 ppdiblcb = -1.028565910e-12
+ drout = 2.747894712e+00 ldrout = -8.685602921e-07 wdrout = -2.592964732e-06 pdrout = 1.267622668e-12
+ pscbe1 = 7.837979489e+08 lpscbe1 = 3.645196149e+00 wpscbe1 = -1.552976458e+00 ppscbe1 = 7.592036010e-7
+ pscbe2 = 1.025310421e-08 lpscbe2 = -4.964784350e-16 wpscbe2 = -1.888406470e-15 ppscbe2 = 9.231852710e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.100425080e+01 lbeta0 = -8.420291984e-07 wbeta0 = -2.419108794e-06 pbeta0 = 1.182629716e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.236382180e-09 lagidl = -5.555431564e-16 wagidl = -2.324608388e-15 pagidl = 1.136431303e-21
+ bgidl = 1.139174799e+09 lbgidl = 2.760937388e+01 wbgidl = 4.200444459e+02 pbgidl = -2.053471283e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.325917527e-01 lkt1 = 6.901463475e-08 wkt1 = 2.839386528e-07 pkt1 = -1.388090892e-13
+ kt2 = -3.966831155e-02 lkt2 = -3.878053400e-09 wkt2 = -1.172510494e-08 pkt2 = 5.732052052e-15
+ at = -1.486758419e+05 lat = 8.979360882e-02 wat = 3.583886969e-01 pat = -1.752054822e-7
+ ute = -1.421594275e-01 lute = 5.972007931e-08 wute = 2.108009942e-07 pute = -1.030542820e-13
+ ua1 = -2.270113440e-09 lua1 = 2.161496388e-15 wua1 = 9.769695213e-15 pua1 = -4.776110899e-21
+ ub1 = 3.129669595e-18 lub1 = -2.348174407e-24 wub1 = -1.027452152e-23 pub1 = 5.022905337e-30
+ uc1 = 4.442561789e-10 luc1 = -2.515178360e-16 wuc1 = -9.603113940e-16 puc1 = 4.694674312e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 9.663038917e-01 lvth0 = -3.553798034e-07 wvth0 = -3.631498828e-06 pvth0 = 6.132512072e-13
+ k1 = -5.278822047e+00 lk1 = 1.053791069e-06 wk1 = 1.076831321e-05 pk1 = -1.818445051e-12
+ k2 = 1.992327629e+00 lk2 = -3.615543996e-07 wk2 = -3.694594814e-06 pk2 = 6.239062262e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.080150869e+00 ldsub = -8.744890130e-08 wdsub = -8.936089771e-07 pdsub = 1.509037480e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 7.435707193e-01 lvoff = -1.752056084e-07 wvoff = -1.790363311e-06 pvoff = 3.023386523e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.294590018e+00 lnfactor = 6.445678720e-07 wnfactor = 6.586608044e-06 pnfactor = -1.112280500e-12
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 5.437140706e-02 lu0 = -8.488895077e-09 wu0 = -8.674497602e-08 pu0 = 1.464862410e-14
+ ua = 9.752543028e-09 lua = -1.971470892e-15 wua = -2.014575439e-14 pua = 3.402013544e-21
+ ub = -4.117078961e-18 lub = 9.916457734e-25 wub = 1.013327271e-23 pub = -1.711205763e-30
+ uc = -2.527105617e-10 luc = 4.126946513e-17 wuc = 4.217178714e-16 puc = -7.121549695e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.601820286e+05 lvsat = 9.104194187e-02 wvsat = 9.303249708e-01 pvsat = -1.571039778e-7
+ a0 = 1.146392495e+00 la0 = -6.557095375e-08 wa0 = -6.700460731e-07 pa0 = 1.131506804e-13
+ ags = 2.333249928e+01 lags = -3.729071658e-06 wags = -3.810604662e-05 pags = 6.434968093e-12
+ a1 = 0.0
+ a2 = 3.654156037e+00 la2 = -5.051377182e-07 wa2 = -5.161821280e-06 pa2 = 8.716767595e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.292491321e-02 lketa = -2.127372133e-08 wketa = -2.173885329e-07 pketa = 3.671040154e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.361753037e+00 lpclm = 3.540264066e-07 wpclm = 3.617668951e-06 ppclm = -6.109157558e-13
+ pdiblc1 = -1.376095058e+00 lpdiblc1 = 3.103208367e-07 wpdiblc1 = 3.171057399e-06 ppdiblc1 = -5.354964629e-13
+ pdiblc2 = -3.076068581e-02 lpdiblc2 = 6.862893847e-09 wpdiblc2 = 7.012945227e-08 ppdiblc2 = -1.184276061e-14
+ pdiblcb = 4.129851026e+00 lpdiblcb = -7.353389020e-07 wpdiblcb = -7.514164664e-06 ppdiblcb = 1.268916987e-12
+ drout = -4.682108439e+00 ldrout = 9.062445604e-07 wdrout = 9.260588328e-06 pdrout = -1.563835551e-12
+ pscbe1 = 7.967858873e+08 lpscbe1 = 5.427673004e-01 wpscbe1 = 5.546344493e+00 ppscbe1 = -9.366111945e-7
+ pscbe2 = 5.411646669e-09 lpscbe2 = 6.600005278e-16 wpscbe2 = 6.744308822e-15 ppscbe2 = -1.138911431e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.939693167e+00 lbeta0 = 8.454816830e-07 wbeta0 = 8.639674263e-06 pbeta0 = -1.458981793e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.490568983e-09 lagidl = 8.124536679e-16 wagidl = 8.302172815e-15 pagidl = -1.401987923e-21
+ bgidl = 1.869343746e+09 lbgidl = -1.468060825e+02 wbgidl = -1.500158735e+03 pbgidl = 2.533318057e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 7.177281692e-02 lkt1 = -9.923693000e-08 wkt1 = -1.014066617e-06 pkt1 = 1.712454296e-13
+ kt2 = -7.305882895e-02 lkt2 = 4.097939491e-09 wkt2 = 4.187537479e-08 pkt2 = -7.071494540e-15
+ at = 7.516085239e+05 lat = -1.252573176e-01 wat = -1.279959632e+00 pat = 2.161467830e-7
+ ute = 4.162836676e-01 lute = -7.367522280e-08 wute = -7.528606936e-07 pute = 1.271355853e-13
+ ua1 = 2.107320144e-08 lua1 = -3.414521237e-15 wua1 = -3.489176862e-14 pua1 = 5.892172967e-21
+ ub1 = -2.173378374e-17 lub1 = 3.590958692e-24 wub1 = 3.669471972e-23 pub1 = -6.196637320e-30
+ uc1 = -2.013766689e-09 luc1 = 3.356300865e-16 wuc1 = 3.429683550e-15 puc1 = -5.791706611e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.081713941e+00 lvth0 = -1.049051290e-08 wvth0 = 5.181396286e-08 pvth0 = -9.630661277e-15
+ k1 = 4.071238096e-01 lk1 = 1.030285673e-07 wk1 = -1.856282002e-07 pk1 = 3.450271357e-14
+ k2 = 1.863348031e-01 lk2 = -6.227188854e-08 wk2 = -3.889440320e-08 pk2 = 7.229302723e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.081497471e+00 ldsub = -2.823726010e-07 wdsub = -2.328098911e-07 pdsub = 4.327237445e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -4.484278162e-01 lvoff = 2.871335909e-08 wvoff = 9.848429104e-07 pvoff = -1.830527518e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.230554396e+01 lnfactor = -1.818400929e-06 wnfactor = -2.673135008e-05 pnfactor = 4.968556040e-12
+ eta0 = -5.351278317e-03 leta0 = 9.207094210e-08 weta0 = 3.883159789e-06 peta0 = -7.217629099e-13
+ etab = -1.261599351e+00 letab = 2.343773026e-07 wetab = 2.577547717e-06 petab = -4.790887941e-13
+ u0 = 1.705850645e-02 lu0 = -2.408116126e-09 wu0 = -1.859560682e-08 pu0 = 3.456365439e-15
+ ua = 4.099998028e-09 lua = -1.119298659e-15 wua = -9.748913973e-15 pua = 1.812030640e-21
+ ub = -1.495708114e-18 lub = 6.042397150e-25 wub = 5.376526352e-24 pub = -9.993349530e-31
+ uc = -5.736685821e-11 luc = 9.115493085e-18 wuc = 1.160732617e-16 puc = -2.157453716e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.023056426e+05 lvsat = -7.869052632e-02 wvsat = -5.958956974e-01 pvsat = 1.107591333e-7
+ a0 = -6.898956592e+00 la0 = 1.423217109e-06 wa0 = 1.415145174e-05 pa0 = -2.630330335e-12
+ ags = 1.249999831e+00 lags = 2.634467666e-14
+ a1 = 0.0
+ a2 = -1.595100384e+00 la2 = 4.196897862e-07 wa2 = 3.575474744e-06 pa2 = -6.645734907e-13
+ b0 = 5.904230970e-23 lb0 = -1.097419410e-29 wb0 = -1.207782477e-28 pb0 = 2.244905289e-35
+ b1 = 0.0
+ keta = -5.965750302e-01 lketa = 9.730722563e-08 wketa = 4.075606500e-07 pketa = -7.575329802e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.349047126e+00 lpclm = -3.000604809e-07 wpclm = -2.175207151e-06 ppclm = 4.043057532e-13
+ pdiblc1 = 2.189823244e+00 lpdiblc1 = -3.212366621e-07 wpdiblc1 = -3.333371279e-07 ppdiblc1 = 6.195737197e-14
+ pdiblc2 = 5.719952706e-02 lpdiblc2 = -8.795389203e-09 wpdiblc2 = -2.902534233e-08 ppdiblc2 = 5.394940379e-15
+ pdiblcb = 3.433942151e+01 lpdiblcb = -6.424417713e-06 wpdiblcb = -6.098588770e-05 ppdiblcb = 1.133544695e-11
+ drout = -9.552668171e-01 ldrout = 3.047673812e-07 wdrout = -3.311541533e-12 pdrout = 6.155162247e-19
+ pscbe1 = 7.895341633e+08 lpscbe1 = 1.945285156e+00 wpscbe1 = 2.140915229e+01 ppscbe1 = -3.979319137e-6
+ pscbe2 = -3.358980641e-08 lpscbe2 = 7.975642307e-15 wpscbe2 = 8.798849792e-14 ppscbe2 = -1.635442211e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.969833793e+01 lbeta0 = -1.998463693e-06 wbeta0 = -1.235519942e-05 pbeta0 = 2.296460916e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.642108846e-08 lagidl = -2.992607077e-15 wagidl = -3.092114238e-14 pagidl = 5.747312734e-21
+ bgidl = 9.999998475e+08 lbgidl = 2.376335716e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.670853509e-01 lkt1 = 9.517539882e-09 wkt1 = 3.438852216e-07 pkt1 = -6.391794613e-14
+ kt2 = -2.619595634e-02 lkt2 = -4.199926541e-09 wkt2 = -1.487305687e-13 pkt2 = 2.764455076e-20
+ at = 1.811172815e+05 lat = -3.182965858e-02 wat = -4.694036583e-01 pat = 8.724805796e-8
+ ute = 1.325677166e+00 lute = -2.501210147e-07 wute = 8.724083407e-13 pute = -1.621545381e-19
+ ua1 = 4.796705996e-09 lua1 = -7.329459926e-16 wua1 = -3.438854770e-15 pua1 = 6.391799362e-22
+ ub1 = -2.170212456e-18 lub1 = 3.161764694e-25 wub1 = 1.522202020e-30 pub1 = -2.829316898e-37
+ uc1 = -7.606959999e-10 luc1 = 1.365094343e-16 wuc1 = 1.501632464e-15 puc1 = -2.791084260e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.101366082e+00 lvth0 = 2.545798937e-7
+ k1 = 4.212606180e-01 lk1 = 1.291674424e-6
+ k2 = 3.716651602e-02 lk2 = -5.420869610e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.367447726e-01 lvoff = -1.216751986e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.592519036e+00 lnfactor = -9.408788196e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.447690685e-02 lu0 = -2.873188681e-8
+ ua = -6.324241445e-10 lua = 4.503683210e-16
+ ub = 1.868978521e-18 lub = -4.055915651e-24
+ uc = -7.214960068e-11 luc = -7.406433888e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.622213786e+00 la0 = -5.637233290e-8
+ ags = 4.822764082e-01 lags = -4.567173287e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.480298045e-02 lketa = 4.710778082e-07 wketa = 8.881784197e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.042722157e-01 lpclm = -2.880916892e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.362535913e-04 lpdiblc2 = 3.013041483e-9
+ pdiblcb = -3.448804924e-03 lpdiblcb = 3.834829377e-8
+ drout = 0.56
+ pscbe1 = 7.008738872e+08 lpscbe1 = 1.786719392e+3
+ pscbe2 = 9.665980000e-09 lpscbe2 = -6.105490408e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.681322036e-10 lalpha0 = -9.357433760e-15
+ alpha1 = -2.464203913e-11 lalpha1 = 2.491453517e-15 walpha1 = 1.227846222e-31 palpha1 = 2.584939414e-35
+ beta0 = 3.268447993e+00 lbeta0 = -5.365972042e-06 wbeta0 = -5.684341886e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.852343277e-11 lagidl = 1.147528989e-15
+ bgidl = 1.562948962e+09 lbgidl = -1.125271361e+4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.257308181e-01 lkt1 = -5.958518612e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.559870728e-01 lute = 5.256487698e-7
+ ua1 = 2.139764998e-09 lua1 = 7.182700633e-15
+ ub1 = -7.306057684e-19 lub1 = -1.899330897e-23
+ uc1 = 4.338507642e-11 luc1 = 7.645641303e-15 puc1 = 5.293955920e-35
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.08863
+ k1 = 0.4858803
+ k2 = 0.010047076
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.24283192
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.5454489
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0130395126
+ ua = -6.0989319e-10
+ ub = 1.66606982e-18
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.6193936
+ ags = 0.47999155
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.093872372e+00 lvth0 = 4.188063158e-8
+ k1 = 4.522972755e-01 lk1 = 2.682904169e-7
+ k2 = 2.243897693e-02 lk2 = -9.899728555e-08 pk2 = 8.881784197e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.402497948e-01 lvoff = -2.062826246e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.707115507e+00 lnfactor = -1.291533511e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.609958679e-02 lu0 = -2.444653486e-8
+ ua = -1.211989359e-10 lua = -3.904114865e-15
+ ub = 1.642518584e-18 lub = 1.881477614e-25
+ uc = -1.423307551e-10 luc = 2.646582022e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.212579461e+05 lvsat = -4.868852462e-1
+ a0 = 1.674871402e+00 la0 = -4.432049504e-7
+ ags = 4.562623108e-01 lags = 1.895698069e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.743565127e-02 lketa = 4.952840774e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.109267259e-01 lpclm = 4.562227086e-06 wpclm = -3.552713679e-21 ppclm = 2.131628207e-26
+ pdiblc1 = 0.39
+ pdiblc2 = 3.587787891e-04 lpdiblc2 = -5.735148984e-10
+ pdiblcb = -4.459427061e-04 lpdiblcb = -8.662970003e-9
+ drout = 0.56
+ pscbe1 = 7.805463027e+08 lpscbe1 = 7.759826970e+1
+ pscbe2 = 9.153007757e-09 lpscbe2 = 1.657912159e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.819567689e-01 lbeta0 = 2.941467397e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.917358547e-10 lagidl = -3.659223987e-16
+ bgidl = 8.022575536e+08 lbgidl = 1.579738698e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.101376581e-01 lkt1 = 4.361735931e-7
+ kt2 = -3.138933667e-02 lkt2 = -5.250016399e-8
+ at = -1.789107917e+05 lat = 1.429295056e+0
+ ute = 1.617288118e-01 lute = -3.925881003e-6
+ ua1 = 5.328096354e-09 lua1 = -2.260048410e-14
+ ub1 = -4.224512371e-18 lub1 = 2.032138745e-23
+ uc1 = 7.901037197e-10 luc1 = -2.909735948e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.091123626e+00 lvth0 = 3.091624109e-8
+ k1 = 5.977558582e-01 lk1 = -3.119249599e-7
+ k2 = -2.975396524e-02 lk2 = 1.091935757e-07 wk2 = -2.220446049e-22 pk2 = 5.551115123e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.223229514e-01 lvoff = -9.213611045e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.717805832e+00 lnfactor = -1.334175826e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.150387845e-03 lu0 = 7.261786318e-9
+ ua = -1.665485757e-09 lua = 2.255844507e-15
+ ub = 2.098150966e-18 lub = -1.629310578e-24
+ uc = -6.694967090e-11 luc = -3.602714318e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.447013512e+05 lvsat = -1.815109412e-1
+ a0 = 1.964115559e+00 la0 = -1.596962289e-6
+ ags = 6.423764338e-01 lags = -5.528152347e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.118284482e-02 lketa = 6.447547569e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.336218480e-01 lpclm = -1.199889384e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 1.963998626e-02 lpdiblcb = -8.878312947e-08 wpdiblcb = -1.110223025e-22 ppdiblcb = -6.661338148e-28
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.671893803e-08 lpscbe2 = -2.852160011e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.565947440e+00 lbeta0 = 4.492596311e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.143013757e+09 lbgidl = 2.205064997e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.434839429e-01 lkt1 = -2.285864121e-7
+ kt2 = -4.017360155e-02 lkt2 = -1.746087337e-8
+ at = 2.745973838e+05 lat = -3.796900997e-1
+ ute = -1.640382899e+00 lute = 3.262508336e-6
+ ua1 = -3.274541222e-09 lua1 = 1.171431885e-14 wua1 = 2.646977960e-29 pua1 = 2.646977960e-35
+ ub1 = 3.170152177e-18 lub1 = -9.174968124e-24 wub1 = 2.465190329e-38 pub1 = -9.860761315e-44
+ uc1 = 9.216446460e-11 luc1 = -1.257469911e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.090838253e+00 lvth0 = 3.034867045e-8
+ k1 = 4.322967437e-01 lk1 = 1.715170913e-8
+ k2 = 2.844424485e-02 lk2 = -6.555098444e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.916658762e-01 ldsub = 3.347946888e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.996927125e-01 lvoff = 6.174228629e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.177495674e-01 lnfactor = 1.649241077e-6
+ eta0 = -5.744849986e-02 leta0 = 2.733671979e-7
+ etab = 6.842919891e-01 letab = -1.500188708e-06 wetab = 5.329070518e-21 petab = -1.776356839e-27
+ u0 = 1.359283912e-02 lu0 = -3.562541745e-9
+ ua = -1.917591780e-10 lua = -6.752060745e-16
+ ub = 1.151418582e-18 lub = 2.536170597e-25
+ uc = -1.214437714e-10 luc = 7.235453841e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.038194939e+04 lvsat = 2.596678738e-2
+ a0 = 1.115812466e+00 la0 = 9.020228253e-8
+ ags = 1.549979248e-01 lags = 4.165172605e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.629453859e-03 lketa = -1.220220699e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.108255342e-02 lpclm = 5.752552428e-7
+ pdiblc1 = 4.088045794e-01 lpdiblc1 = -3.739986375e-8
+ pdiblc2 = 2.392950000e-06 lpdiblc2 = 4.228477835e-10
+ pdiblcb = -0.025
+ drout = 1.344068365e-01 ldrout = 8.464494752e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.454152232e-09 lpscbe2 = 1.358892391e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.794355910e+00 lbeta0 = 2.049451557e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.269088568e+09 lbgidl = -3.023991007e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444605805e-01 lkt1 = -2.775700689e-8
+ kt2 = -6.040588351e-02 lkt2 = 2.277850526e-8
+ at = 6.493100483e+04 lat = 3.730907145e-2
+ ute = 0.0
+ ua1 = 2.824339679e-09 lua1 = -4.155624112e-16
+ ub1 = -1.527062104e-18 lub1 = 1.671804431e-25
+ uc1 = 1.528486051e-10 luc1 = -2.464398577e-16 wuc1 = 8.271806126e-31 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.083811263e+00 lvth0 = 2.339989136e-8
+ k1 = 3.328536151e-01 lk1 = 1.154880357e-7
+ k2 = 6.118412774e-02 lk2 = -3.893058644e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.664626476e-01 ldsub = 2.608304055e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.329295969e-01 lvoff = -4.277755777e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.557974615e+00 lnfactor = 3.239327345e-7
+ eta0 = 3.582529886e-01 leta0 = -1.377075330e-7
+ etab = -1.646537114e+00 letab = 8.046982669e-7
+ u0 = 1.168706777e-02 lu0 = -1.677981632e-09 wu0 = 2.220446049e-22
+ ua = -5.906662208e-10 lua = -2.807388671e-16
+ ub = 1.291920204e-18 lub = 1.146792206e-25
+ uc = -6.422249855e-11 luc = 1.577013837e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.500133002e+04 lvsat = 1.621420453e-3
+ a0 = 1.232969442e+00 la0 = -2.565073621e-8
+ ags = -8.543032923e-02 lags = 6.542695481e-7
+ a1 = 0.0
+ a2 = 6.044617774e-01 la2 = 1.933618822e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.631183582e-02 lketa = -3.093268012e-08 pketa = 2.220446049e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.378830106e-01 lpclm = 8.398417474e-8
+ pdiblc1 = -2.440305587e-01 lpdiblc1 = 6.081692192e-7
+ pdiblc2 = -1.444786656e-04 lpdiblc2 = 5.680847180e-10
+ pdiblcb = -4.911716338e-02 lpdiblcb = 2.384873935e-8
+ drout = 1.009114736e+00 ldrout = -1.852292549e-8
+ pscbe1 = 8.085510012e+08 lpscbe1 = -8.455828520e+0
+ pscbe2 = 9.336779542e-09 lpscbe2 = -4.851479500e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.461134792e+00 lbeta0 = 4.012239235e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.280411890e+09 lbgidl = -4.143720287e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.540604914e-01 lkt1 = -1.826394297e-8
+ kt2 = -2.736871980e-02 lkt2 = -9.890954821e-9
+ at = 1.688138884e+05 lat = -6.541759562e-2
+ ute = 1.955480000e-02 lute = -1.933715508e-8
+ ua1 = 2.651272672e-09 lua1 = -2.444216402e-16
+ ub1 = -1.049425256e-18 lub1 = -3.051403071e-25
+ uc1 = -1.219162794e-10 luc1 = 2.526689368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.382883043e-01 lvth0 = -4.774191768e-8
+ k1 = 1.942152608e-01 lk1 = 1.832641680e-7
+ k2 = 1.059965720e-01 lk2 = -6.083804605e-08 pk2 = -4.440892099e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.418210343e+00 ldsub = -2.044504902e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.917397620e-01 lvoff = -2.441423037e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.932257307e+00 lnfactor = 1.409571549e-7
+ eta0 = -3.184587778e-01 leta0 = 1.931165483e-07 weta0 = -1.776356839e-21
+ etab = -3.801533128e-04 letab = -5.848652817e-11
+ u0 = 1.222195773e-02 lu0 = -1.939473286e-09 wu0 = -2.220446049e-22
+ ua = -4.416108828e-10 lua = -3.536075502e-16
+ ub = 1.308016311e-18 lub = 1.068103164e-25
+ uc = -5.455131315e-11 luc = 1.104218596e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.816660043e+04 lvsat = 4.962714709e-3
+ a0 = 1.584094753e+00 la0 = -1.973053668e-7
+ ags = 1.255670918e+00 lags = -1.354618715e-9
+ a1 = 0.0
+ a2 = 1.322097146e+00 la2 = -1.574685206e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.203352684e-02 lketa = -1.218678267e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.857741658e-01 lpclm = 1.168462571e-8
+ pdiblc1 = 1.514491131e+00 lpdiblc1 = -2.515192790e-07 wpdiblc1 = -2.842170943e-20
+ pdiblc2 = -7.449769845e-03 lpdiblc2 = 4.139422417e-09 wpdiblc2 = -2.775557562e-23 ppdiblc2 = -2.081668171e-29
+ pdiblcb = 2.139637357e-01 lpdiblcb = -1.047636198e-07 wpdiblcb = -2.359223927e-22 ppdiblcb = -4.475586568e-28
+ drout = 1.245268568e+00 ldrout = -1.339714492e-7
+ pscbe1 = 7.828979972e+08 lpscbe1 = 4.085155538e+0
+ pscbe2 = 9.158770415e-09 lpscbe2 = 3.850852687e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.602374377e+00 lbeta0 = -1.566938724e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.107311437e-10 lagidl = 1.030201342e-16 pagidl = 8.271806126e-37
+ bgidl = 1.382591054e+09 lbgidl = -9.138953103e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.680489659e-01 lkt1 = -1.142539742e-8
+ kt2 = -4.646302380e-02 lkt2 = -5.563224232e-10
+ at = 5.901083391e+04 lat = -1.173817637e-2
+ ute = -2.000000080e-02 lute = 3.899890411e-16
+ ua1 = 3.391436548e-09 lua1 = -6.062655543e-16
+ ub1 = -2.824427839e-18 lub1 = 5.626052055e-25
+ uc1 = -1.122454153e-10 luc1 = 2.053909835e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.13815399562893
+ k1 = 0.961428255393082
+ k2 = -0.148694456831761
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.562303405039308
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.293946947389937
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.5223571722327
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 0.0041025903490566
+ ua = -1.92194558459119e-9
+ ub = 1.75516461966667e-18
+ uc = -8.324553995283e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 78942.397761062
+ a0 = 0.758099999261006
+ ags = 1.24999997272013
+ a1 = 0.0
+ a2 = 0.662874470440252
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0730519999606918
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.734690420259434
+ pdiblc1 = 0.461536473183962
+ pdiblc2 = 0.00987941513820755
+ pdiblcb = -0.224616327814465
+ drout = 0.684413503600629
+ pscbe1 = 800000000.518868
+ pscbe2 = 9.31998164677673e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.94639467130503
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.20550031084906e-10
+ bgidl = 999999975.393082
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.515879992940252
+ kt2 = -0.0487919994941038
+ at = 9870.39612421382
+ ute = -0.0199999991650943
+ ua1 = 8.53380055896226e-10
+ ub1 = -4.69150049528303e-19
+ uc1 = -2.62609955581761e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.051692103e+00 lvth0 = -1.607067203e-08 wvth0 = 7.617756864e-12 pvth0 = -1.415912479e-18
+ k1 = 2.995547351e-01 lk1 = 1.230224312e-07 wk1 = -4.638744258e-12 pk1 = 8.622033931e-19
+ k2 = 1.637940389e-01 lk2 = -5.808223670e-08 wk2 = 2.435342125e-12 pk2 = -4.526570372e-19
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.946566500e+00 ldsub = -2.572929815e-07 wdsub = 2.996034488e-11 pdsub = -5.568729293e-18
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.222785319e-01 lvoff = -7.736382983e-08 wvoff = 1.948060753e-11 pvoff = -3.620860525e-18
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -3.185176667e+00 lnfactor = 1.060859315e-06 wnfactor = -2.217650692e-10 pnfactor = 4.121947342e-17
+ eta0 = 2.244936646e+00 leta0 = -3.261900743e-07 weta0 = 1.344066141e-11 peta0 = -2.498215743e-18
+ etab = 2.320943525e-01 letab = -4.325554605e-08 wetab = -2.999119890e-12 petab = 5.574464145e-19
+ u0 = 6.282310451e-03 lu0 = -4.051445754e-10 wu0 = 3.407776283e-14 pu0 = -6.334033797e-21
+ ua = -1.549498325e-09 lua = -6.922677217e-17 wua = -1.877841360e-20 pua = 3.490343731e-27
+ ub = 1.620010242e-18 lub = 2.512114415e-26 wub = -2.578973141e-29 pub = 4.793537375e-36
+ uc = 9.897706192e-12 luc = -3.386971501e-18 wuc = 4.957926535e-23 puc = -9.215298052e-30
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.569838217e+05 lvsat = -1.450555947e-02 wvsat = -7.661910579e-07 pvsat = 1.424119323e-13
+ a0 = 1.301824142e+00 la0 = -1.010620064e-07 wa0 = 4.089757397e-12 pa0 = -7.601632177e-19
+ ags = 1.249999831e+00 lags = 2.634469354e-14
+ a1 = 0.0
+ a2 = 4.768820509e-01 la2 = 3.457041102e-08 wa2 = 1.627072265e-11 pa2 = -3.024239220e-18
+ b0 = -1.094875900e-23 lb0 = 2.035045836e-30 wb0 = -1.196924258e-34 pb0 = 2.224723122e-41
+ b1 = 0.0
+ keta = -3.603916731e-01 lketa = 5.340782504e-08 wketa = -2.547054891e-12 pketa = 4.734210934e-19
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.088513738e+00 lpclm = -6.576514013e-08 wpclm = -3.005929216e-12 ppclm = 5.587120597e-19
+ pdiblc1 = 1.996662586e+00 lpdiblc1 = -2.853338906e-07 wpdiblc1 = -1.484718064e-11 ppdiblc1 = 2.759645469e-18
+ pdiblc2 = 4.037920184e-02 lpdiblc2 = -5.668995354e-09 wpdiblc2 = 1.809217531e-13 ppdiblc2 = -3.362792622e-20
+ pdiblcb = -1.001973283e+00 lpdiblcb = 1.444873373e-07 wpdiblcb = 6.702776716e-13 ppdiblcb = -1.245845063e-19
+ drout = -9.552857037e-01 ldrout = 3.047708917e-07 wdrout = 2.927942791e-11 pdrout = -5.442167264e-18
+ pscbe1 = 8.019400484e+08 lpscbe1 = -3.605966932e-01 wpscbe1 = 1.284166687e-03 ppscbe1 = -2.386880646e-10
+ pscbe2 = 1.739956503e-08 lpscbe2 = -1.501752163e-15 wpscbe2 = 1.167985276e-19 ppscbe2 = -2.170934231e-26
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.253849864e+01 lbeta0 = -6.676643648e-07 wbeta0 = -2.323415902e-11 pbeta0 = 4.318533342e-18
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.497745042e-09 lagidl = 3.379665052e-16 wagidl = -9.082793639e-21 pagidl = 1.688218853e-27
+ bgidl = 9.999998475e+08 lbgidl = 2.376335144e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.678029168e-01 lkt1 = -2.752308615e-08 wkt1 = -9.309413258e-13 pkt1 = 1.730340671e-19
+ kt2 = -2.619680459e-02 lkt2 = -4.199768877e-09 wkt2 = 1.315020793e-12 pkt2 = -2.444229148e-19
+ at = -9.090145530e+04 lat = 1.873046402e-02 wat = -2.141696499e-06 pat = 3.980771280e-13
+ ute = 1.325682142e+00 lute = -2.501219395e-07 wute = -7.713512574e-12 pute = 1.433710575e-18
+ ua1 = 2.803882499e-09 lua1 = -3.625398891e-16 wua1 = 5.298384738e-21 pua1 = -9.848107706e-28
+ ub1 = -2.170203774e-18 lub1 = 3.161748558e-25 wub1 = -1.345874841e-29 pub1 = 2.501577567e-36
+ uc1 = 1.095003338e-10 luc1 = -2.523395829e-17 wuc1 = 2.525776211e-21 puc1 = -4.694660250e-28
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.121519770e+00 lvth0 = -1.141251892e-06 wvth0 = 3.417303649e-08 pvth0 = 2.366803085e-12
+ k1 = 1.728409333e-01 lk1 = 8.824441367e-06 wk1 = 4.212258826e-07 pk1 = -1.277272535e-11
+ k2 = 1.375340493e-01 lk2 = -3.314597553e-06 wk2 = -1.701853975e-07 pk2 = 4.701129955e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.082678163e-01 lvoff = -1.338794682e-06 wvoff = -4.828615362e-08 pvoff = 2.063774574e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.249600278e+00 lnfactor = -5.403537089e-05 wnfactor = -1.114161411e-06 pnfactor = 9.002818884e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.638637523e-02 lu0 = 1.653053085e-07 wu0 = -3.237736590e-09 pu0 = -3.290137371e-13
+ ua = -7.471786972e-10 lua = 5.890308438e-15 wua = 1.945803441e-16 pua = -9.224082141e-21
+ ub = 2.011695620e-18 lub = 3.601695043e-23 wub = -2.419942532e-25 pub = -6.794843333e-29
+ uc = 8.319917263e-11 luc = -6.350317454e-15 wuc = -2.634127977e-16 puc = 9.511886758e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.603104088e+05 lvsat = 2.090945812e-04 wvsat = 3.545848372e-06 pvsat = -3.545453719e-10
+ a0 = 1.401868330e+00 la0 = 2.273102276e-05 wa0 = 3.736226027e-07 pa0 = -3.863880845e-11
+ ags = 2.146649182e-01 lags = 2.732442923e-05 wags = 4.537679298e-07 pags = -4.640934533e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.091357611e-01 lketa = -4.079618329e-07 wketa = 9.212785820e-08 pketa = 1.490518954e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.543676277e-01 lpclm = -1.928451140e-05 wpclm = -9.327538827e-07 ppclm = 2.781429574e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -3.413474094e-04 lpdiblc2 = 1.039773684e-08 wpdiblc2 = 8.098307639e-10 ppdiblc2 = -1.252165192e-14
+ pdiblcb = -1.383443847e-01 lpdiblcb = 1.301259714e-05 wpdiblcb = 2.287319127e-07 ppdiblcb = -2.199942178e-11
+ drout = 0.56
+ pscbe1 = 4.097397702e+08 lpscbe1 = 6.957618348e+03 wpscbe1 = 4.936534138e+02 ppscbe1 = -8.767890029e-3
+ pscbe2 = 7.396955570e-09 lpscbe2 = 3.025758131e-13 wpscbe2 = 3.847407743e-15 ppscbe2 = -5.234068093e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.135321188e-09 lalpha0 = -4.068377063e-14 walpha0 = -2.657360120e-15 palpha0 = 5.311762598e-20
+ alpha1 = -4.419122658e-10 lalpha1 = 1.083221383e-14 walpha1 = 7.075325764e-16 palpha1 = -1.414277669e-20
+ beta0 = 6.909590680e+00 lbeta0 = -2.975440007e-04 wbeta0 = -6.174001644e-06 pbeta0 = 4.954234933e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.465782709e-10 lagidl = -2.003241973e-14 wagidl = -9.843906074e-17 pagidl = 3.591318701e-20
+ bgidl = 3.447560627e+09 lbgidl = -4.892397119e+04 wbgidl = -3.195589001e+03 pbgidl = 6.387621311e-2
+ cgidl = 300.0
+ egidl = 7.570061872e-01 legidl = -6.569330624e-05 wegidl = -1.114034145e-06 pegidl = 1.113910153e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.135837395e-01 lkt1 = -3.825819494e-06 wkt1 = -1.901590537e-07 pkt1 = 5.476804178e-12
+ kt2 = -5.000407391e-02 lkt2 = 1.204173351e-06 wkt2 = 2.042050106e-08 pkt2 = -2.041822826e-12
+ at = 0.0
+ ute = -2.788836306e-01 lute = -1.422671664e-05 wute = -1.307382929e-07 pute = 2.501443533e-11
+ ua1 = 3.710327627e-10 lua1 = 8.779917495e-14 wua1 = 2.999101291e-15 pua1 = -1.366950674e-19
+ ub1 = 3.257526331e-18 lub1 = -1.632812093e-22 wub1 = -6.762364526e-24 pub1 = 2.446577382e-28
+ uc1 = -1.600676817e-09 luc1 = 6.959378104e-14 wuc1 = 2.787707516e-15 puc1 = -1.050406286e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.178614138e+00 wvth0 = 1.525790837e-7
+ k1 = 6.143086784e-01 wk1 = -2.177659839e-7
+ k2 = -2.828810839e-02 wk2 = 6.500198203e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.752448231e-01 wvoff = 5.496003156e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -4.536726379e-01 wnfactor = 3.389754460e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.465624283e-02 wu0 = -1.969758335e-8
+ ua = -4.524992862e-10 wua = -2.668805660e-16
+ ub = 3.813545872e-18 wub = -3.641307637e-24
+ uc = -2.344934960e-10 wuc = 2.124463558e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.603208694e+05 wvsat = -1.419129094e-5
+ a0 = 2.539052311e+00 wa0 = -1.559393543e-6
+ ags = 1.581647105e+00 wags = -1.867991396e-6
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.295452106e-01 wketa = 1.666953027e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.103948328e-01 wpclm = 4.587352678e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.788289110e-04 wpdiblc2 = 1.833995591e-10
+ pdiblcb = 5.126477496e-01 wpdiblcb = -8.718516511e-7
+ drout = 0.56
+ pscbe1 = 7.578143911e+08 wpscbe1 = 5.501480994e+1
+ pscbe2 = 2.253417009e-08 wpscbe2 = -2.233750462e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -7.975893126e+00 wbeta0 = 1.861096585e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.556004282e-10 wagidl = 1.698220131e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -2.529488059e+00 wegidl = 4.458617801e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.049812269e-01 wkt1 = 8.383363211e-8
+ kt2 = 1.023811843e-02 wkt2 = -8.172748559e-8
+ at = 0.0
+ ute = -9.906155412e-01 wute = 1.120679888e-6
+ ua1 = 4.763435883e-09 wua1 = -3.839457738e-15
+ ub1 = -4.911079965e-18 wub1 = 5.477333775e-24
+ uc1 = 1.880949760e-09 wuc1 = -2.467248297e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.180788490e+00 lvth0 = 1.737061476e-08 wvth0 = 1.473768807e-07 pvth0 = 4.155972373e-14
+ k1 = 4.412317095e-01 lk1 = 1.382689405e-06 wk1 = 1.876301716e-08 pk1 = -1.889599441e-12
+ k2 = 3.434970078e-02 lk2 = -5.004053146e-07 wk2 = -2.019608540e-08 pk2 = 6.806362850e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.914841189e-01 lvoff = 1.297336230e-07 wvoff = 8.687404706e-08 pvoff = -2.549569210e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.436458128e+00 lnfactor = 7.851345515e-06 wnfactor = 5.330312614e-06 pnfactor = -1.550286682e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.905935495e-02 lu0 = -1.150645903e-07 wu0 = -3.893108801e-08 pu0 = 1.536539684e-13
+ ua = 1.800356156e-09 lua = -1.799776925e-14 wua = -3.258231087e-15 pua = 2.389751044e-20
+ ub = 3.684350605e-18 lub = 1.032124187e-24 wub = -3.462175295e-24 pub = -1.431064994e-30
+ uc = -3.816433969e-10 luc = 1.175561429e-15 wuc = 4.057837803e-16 puc = -1.544547551e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.851127815e+04 lvsat = 7.334548890e-01 wvsat = 2.590006106e-01 pvsat = -2.069235581e-6
+ a0 = 2.669974039e+00 la0 = -1.045916665e-06 wa0 = -1.687317923e-06 pa0 = 1.021971243e-12
+ ags = 1.685678218e+00 lags = -8.310910352e-07 wags = -2.084624659e-06 pags = 1.730654978e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.599307534e-01 lketa = 2.427461510e-07 wketa = 2.077053900e-07 pketa = -3.276242562e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.024352626e+00 lpclm = 2.248034299e-05 wpclm = 4.261820251e-06 ppclm = -3.038235153e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 6.189427901e-03 lpdiblc2 = -4.801789395e-08 wpdiblc2 = -9.886576909e-09 ppdiblc2 = 8.044773290e-14
+ pdiblcb = 8.302761565e-01 lpdiblcb = -2.537492052e-06 wpdiblcb = -1.408590667e-06 ppdiblcb = 4.287938225e-12
+ drout = 0.56
+ pscbe1 = -7.024619961e+08 lpscbe1 = 1.166595822e+04 wpscbe1 = 2.514621498e+03 ppscbe1 = -1.964947808e-2
+ pscbe2 = 9.644516451e-08 lpscbe2 = -5.904653260e-13 wpscbe2 = -1.480145014e-13 ppscbe2 = 1.004017189e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.452847448e+01 lbeta0 = 5.234772057e-05 wbeta0 = 2.347846005e-05 pbeta0 = -3.888577834e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.475712186e-09 lagidl = 4.953992219e-15 wagidl = 2.827361582e-15 pagidl = -9.020564264e-21
+ bgidl = 1.402655322e+08 lbgidl = 6.868306898e+03 wbgidl = 1.122488235e+03 pbgidl = -8.967412588e-3
+ cgidl = 300.0
+ egidl = -5.151659567e+00 legidl = 2.094818730e-05 wegidl = 8.904829498e-06 pegidl = -3.552020724e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.573955395e-01 lkt1 = 2.815392129e-06 wkt1 = 5.888181033e-07 pkt1 = -4.034255293e-12
+ kt2 = 2.564819125e-02 lkt2 = -1.231090685e-07 wkt2 = -9.671408718e-08 pkt2 = 1.197260119e-13
+ at = -4.751433594e+05 lat = 3.795858529e+00 wat = 5.022984589e-01 pat = -4.012797089e-6
+ ute = 1.253668267e+00 lute = -1.792929159e-05 wute = -1.851516563e-06 pute = 2.374449106e-11
+ ua1 = 2.121980371e-08 lua1 = -1.314677833e-13 wua1 = -2.694632861e-14 pua1 = 1.845977875e-19
+ ub1 = -2.108101345e-17 lub1 = 1.291794966e-22 wub1 = 2.858225408e-23 pub1 = -1.845822047e-28
+ uc1 = 3.474085516e-09 luc1 = -1.272735444e-14 wuc1 = -4.551018581e-15 puc1 = 1.664696991e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.201895256e+00 lvth0 = 1.015627603e-07 wvth0 = 1.878268116e-07 pvth0 = -1.197897921e-13
+ k1 = 1.116679585e+00 lk1 = -1.311584361e-06 wk1 = -8.798984869e-07 pk1 = 1.695044473e-12
+ k2 = -2.021138318e-01 lk2 = 4.428169765e-07 wk2 = 2.922571816e-07 pk2 = -5.656991782e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.344110573e-01 ldsub = 3.966576434e-06 wdsub = 1.686145266e-06 pdsub = -6.725814266e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -7.812428744e-02 lvoff = -7.213310078e-07 wvoff = -2.445064269e-07 pvoff = 1.066876710e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 4.670774756e+00 lnfactor = -1.650961252e-05 wnfactor = -5.007119073e-06 pnfactor = 2.573180432e-11
+ eta0 = -1.846649205e-01 leta0 = 1.055713961e-06 weta0 = 4.487716618e-07 peta0 = -1.790091818e-12
+ etab = 1.613778929e-01 letab = -9.229363358e-07 wetab = -3.923294456e-07 petab = 1.564951156e-12
+ u0 = 5.689185859e-03 lu0 = 1.804467609e-08 wu0 = 4.173268235e-09 pu0 = -1.828370511e-14
+ ua = -4.699980971e-09 lua = 7.931230499e-15 wua = 5.145356843e-15 pua = -9.623309348e-21
+ ub = 5.742820689e-18 lub = -7.178845374e-24 wub = -6.179982164e-24 pub = 9.409913290e-30
+ uc = -3.814362266e-11 luc = -1.946145158e-16 wuc = -4.884416912e-17 puc = 2.689042380e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.502281180e+05 lvsat = -7.891639620e-01 wvsat = -5.180579075e-01 pvsat = 1.030349830e-6
+ a0 = 4.078328353e+00 la0 = -6.663658935e-06 wa0 = -3.584905726e-06 pa0 = 8.591202300e-12
+ ags = 2.293131095e+00 lags = -3.254141592e-06 wags = -2.799055920e-06 pags = 4.580428401e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.005320765e-01 lketa = 4.046995508e-07 wketa = 2.701960629e-07 pketa = -5.768914267e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.886142155e+00 lpclm = -1.306246232e-05 wpclm = -8.397602387e-06 ppclm = 2.011443965e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.116257839e-02 lpdiblc2 = 2.119700338e-08 wpdiblc2 = 1.929207222e-08 ppdiblc2 = -3.594210526e-14
+ pdiblcb = 4.120466754e-01 lpdiblcb = -8.692290214e-07 wpdiblcb = -6.653734151e-07 ppdiblcb = 1.323341224e-12
+ drout = 0.56
+ pscbe1 = 3.610583925e+09 lpscbe1 = -5.538221261e+03 wpscbe1 = -4.765687936e+03 ppscbe1 = 9.390729811e-3
+ pscbe2 = -8.202937486e-08 lpscbe2 = 1.214464098e-13 wpscbe2 = 1.674398118e-13 ppscbe2 = -2.542890569e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.407591857e+01 lbeta0 = 5.054253387e-05 wbeta0 = 3.330518012e-05 pbeta0 = -7.808328723e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.647896972e-10 lagidl = 9.215538311e-16 wagidl = 9.576698360e-16 pagidl = -1.562606950e-21
+ bgidl = 1.621787880e+09 lbgidl = 9.587068515e+02 wbgidl = -8.118199350e+02 pbgidl = -1.251708757e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.185754887e-01 lkt1 = -1.077629426e-06 wkt1 = -7.834781375e-07 pkt1 = 1.439656013e-12
+ kt2 = 2.693027371e-02 lkt2 = -1.282231287e-07 wkt2 = -1.137828072e-07 pkt2 = 1.878109170e-13
+ at = 8.520883640e+05 lat = -1.498296275e+00 wat = -9.792064107e-01 pat = 1.896733240e-6
+ ute = -6.689477486e+00 lute = 1.375488421e-05 wute = 8.561355863e-06 pute = -1.779110337e-11
+ ua1 = -2.534903998e-08 lua1 = 5.428928029e-14 wua1 = 3.743000574e-14 pua1 = -7.219104127e-20
+ ub1 = 2.326426416e-17 lub1 = -4.770805098e-23 wub1 = -3.407201836e-23 pub1 = 6.533754302e-29
+ uc1 = 3.412091491e-10 luc1 = -2.307178918e-16 wuc1 = -4.222856460e-16 puc1 = 1.779909686e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.152218003e+00 lvth0 = 2.761162340e-09 wvth0 = 1.040768541e-07 pvth0 = 4.677798568e-14
+ k1 = 6.850095563e-01 lk1 = -4.530487916e-07 wk1 = -4.285054047e-07 pk1 = 7.972823134e-13
+ k2 = -6.581041321e-02 lk2 = 1.717271965e-07 wk2 = 1.598202718e-07 pk2 = -3.022993814e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.534590227e+00 ldsub = -1.938381150e-06 wdsub = -3.633589673e-06 pdsub = 3.854446962e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -5.798958062e-01 lvoff = 2.766273127e-07 wvoff = 4.751185302e-07 pvoff = -3.643637783e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -6.756371929e+00 lnfactor = 6.217496709e-06 wnfactor = 1.182547384e-05 pnfactor = -7.746034751e-12
+ eta0 = 4.752066603e-01 leta0 = -2.566848296e-07 weta0 = -9.031818080e-07 peta0 = 8.987678790e-13
+ etab = 2.443710575e-01 letab = -1.087998951e-06 wetab = 7.459396098e-07 petab = -6.989180207e-13
+ u0 = 1.584083623e-02 lu0 = -2.145636793e-09 wu0 = -3.811753363e-09 pu0 = -2.402535207e-15
+ ua = 2.013489644e-10 lua = -1.816877568e-15 wua = -6.665628147e-16 pua = 1.935843302e-21
+ ub = 1.027159610e-18 lub = 2.199991475e-24 wub = 2.106962456e-25 pub = -3.300315278e-30
+ uc = -2.772127238e-10 luc = 2.808628473e-16 wuc = 2.641252626e-16 puc = -3.535512757e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.338136527e+04 lvsat = 1.527837310e-01 wvsat = 1.081184791e-01 pvsat = -2.150335996e-7
+ a0 = 2.399737491e-01 la0 = 9.703293851e-07 wa0 = 1.485091397e-06 pa0 = -1.492362878e-12
+ ags = 2.682639906e-01 lags = 7.730558451e-07 wags = -1.920564330e-07 pags = -6.045546679e-13
+ a1 = 0.0
+ a2 = 1.462064550e+00 la2 = -1.316760322e-06 wa2 = -1.122611217e-06 pa2 = 2.232727770e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.488727691e-02 lketa = -4.363023861e-08 wketa = -4.665797406e-08 pketa = 5.329006183e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.364808545e+00 lpclm = 1.358735996e-06 wpclm = 2.383859876e-06 ppclm = -1.328487202e-12
+ pdiblc1 = -6.902237986e-01 lpdiblc1 = 2.148424706e-06 wpdiblc1 = 1.863536696e-06 ppdiblc1 = -3.706332229e-12
+ pdiblc2 = -1.429128003e-03 lpdiblc2 = 1.838435909e-09 wpdiblc2 = 2.427318422e-09 ppdiblc2 = -2.400302368e-15
+ pdiblcb = -0.025
+ drout = 1.662427097e-01 ldrout = 7.831320619e-07 wdrout = -5.398160712e-08 pdrout = 1.073623989e-13
+ pscbe1 = 8.063185820e+08 lpscbe1 = 3.909795145e+01 wpscbe1 = -1.071392670e+01 ppscbe1 = -6.629534663e-5
+ pscbe2 = -5.125104139e-08 lpscbe2 = 6.023230573e-14 wpscbe2 = 7.934983478e-14 ppscbe2 = -7.908954437e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.811074221e+00 lbeta0 = 3.034410532e-06 wbeta0 = -5.115213936e-06 pbeta0 = -1.670118107e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.249128261e-09 lagidl = -2.487206179e-15 wagidl = -1.948487161e-15 pagidl = 4.217361516e-21
+ bgidl = 2.169929479e+09 lbgidl = -1.314755302e+02 wbgidl = -1.527485666e+03 pbgidl = 1.716573447e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.961606329e-01 lkt1 = -5.388619587e-08 wkt1 = -8.189845366e-08 pkt1 = 4.430522768e-14
+ kt2 = -7.474559650e-02 lkt2 = 7.399695926e-08 wkt2 = 2.431473282e-08 pkt2 = -8.684713741e-14
+ at = -4.051388487e+04 lat = 2.769735598e-01 wat = 1.787946748e-01 pat = -4.063803790e-7
+ ute = -3.019537603e+00 lute = 6.455850877e-06 wute = 5.119994390e-06 pute = -1.094668278e-11
+ ua1 = -7.887599455e-09 lua1 = 1.956074506e-14 wua1 = 1.816339966e-14 pua1 = -3.387226643e-20
+ ub1 = 7.362582748e-18 lub1 = -1.608167386e-23 wub1 = -1.507347738e-23 pub1 = 2.755191483e-29
+ uc1 = 1.083744252e-09 luc1 = -1.707523682e-15 wuc1 = -1.578447138e-15 puc1 = 2.477445876e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.164758661e+00 lvth0 = 1.516224349e-08 wvth0 = 1.372561889e-07 pvth0 = 1.396793696e-14
+ k1 = -2.814058615e-01 lk1 = 5.026104226e-07 wk1 = 1.041551882e-06 pk1 = -6.564132359e-13
+ k2 = 2.783693339e-01 lk2 = -1.686218301e-07 wk2 = -3.682640137e-07 pk2 = 2.199073260e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.255588468e+00 ldsub = 2.798482856e-06 wdsub = 4.615569756e-06 pdsub = -4.302899323e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -3.475471222e-01 lvoff = 4.686466953e-08 wvoff = 1.943479974e-07 pvoff = -8.671822148e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 6.909357503e-01 lnfactor = -1.146922436e-06 wnfactor = 1.470170173e-06 pnfactor = 2.494014386e-12
+ eta0 = 1.704860769e+00 leta0 = -1.472652888e-06 weta0 = -2.283337777e-06 peta0 = 2.263562712e-12
+ etab = -1.692616665e+00 letab = 8.274300984e-07 wetab = 7.813350071e-08 petab = -3.854459355e-14
+ u0 = 2.398927227e-02 lu0 = -1.020338074e-08 wu0 = -2.085988860e-08 pu0 = 1.445585428e-14
+ ua = 2.967851474e-11 lua = -1.647117811e-15 wua = -1.051870181e-15 pua = 2.316862197e-21
+ ub = 3.364902026e-18 lub = -1.117318676e-25 wub = -3.514993583e-24 pub = 3.839076222e-31
+ uc = 5.203953773e-11 luc = -4.472483652e-17 wuc = -1.971364665e-16 puc = 1.025766103e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.150997550e+05 lvsat = 1.584390562e-02 wvsat = -8.494799154e-02 pvsat = -2.411595874e-8
+ a0 = -2.577680633e-01 la0 = 1.462531331e-06 wa0 = 2.527727311e-06 pa0 = -2.523394253e-12
+ ags = 8.421653082e-01 lags = 2.055420491e-07 wags = -1.572851570e-06 pags = 7.608722192e-13
+ a1 = 0.0
+ a2 = -7.520729984e-01 la2 = 8.727338758e-07 wa2 = 2.300170210e-06 pa2 = -1.151958099e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.813442977e-02 lketa = -5.672995066e-08 wketa = -3.700287040e-08 pketa = 4.374241947e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.907425967e+00 lpclm = 2.884184086e-06 wpclm = 5.841941700e-06 ppclm = -4.748080575e-12
+ pdiblc1 = -1.283195189e+00 lpdiblc1 = 2.734796325e-06 wpdiblc1 = 1.762030408e-06 ppdiblc1 = -3.605955706e-12
+ pdiblc2 = -3.343804387e-03 lpdiblc2 = 3.731801944e-09 wpdiblc2 = 5.424847079e-09 ppdiblc2 = -5.364468531e-15
+ pdiblcb = -1.119480211e-01 lpdiblcb = 8.598028965e-08 wpdiblcb = 1.065373847e-07 ppdiblcb = -1.053516236e-13
+ drout = 1.039628582e+00 ldrout = -8.053302554e-08 wdrout = -5.173994838e-08 pdrout = 1.051456899e-13
+ pscbe1 = 9.278700197e+08 lpscbe1 = -8.110061869e+01 wpscbe1 = -2.023199528e+02 ppscbe1 = 1.231781044e-4
+ pscbe2 = 1.036804785e-08 lpscbe2 = -7.009630481e-16 wpscbe2 = -1.748641236e-15 ppscbe2 = 1.106305612e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.466161651e+01 lbeta0 = -1.762145218e-06 wbeta0 = -1.051367321e-05 pbeta0 = 3.668256311e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.298733123e-09 lagidl = 1.021167508e-15 wagidl = 4.067344655e-15 pagidl = -1.731514092e-21
+ bgidl = 2.219160434e+09 lbgidl = -1.801585457e+02 wbgidl = -1.591762685e+03 pbgidl = 2.352189607e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.634902094e-01 lkt1 = 1.115810025e-07 wkt1 = 1.855514374e-07 pkt1 = -2.201679461e-13
+ kt2 = 9.559689512e-02 lkt2 = -9.444962043e-08 wkt2 = -2.085032019e-07 pkt2 = 1.433795337e-13
+ at = 4.398981526e+05 lat = -1.980914917e-01 wat = -4.596564423e-01 pat = 2.249647771e-7
+ ute = 6.374961427e+00 lute = -2.834087378e-06 wute = -1.077636729e-05 pute = 4.772752402e-12
+ ua1 = 2.277750131e-08 lua1 = -1.076305313e-14 wua1 = -3.412647606e-14 pua1 = 1.783562297e-20
+ ub1 = -1.846974694e-17 lub1 = 9.463142001e-24 wub1 = 2.953828070e-23 pub1 = -1.656331438e-29
+ uc1 = -1.612488626e-09 luc1 = 9.587001245e-16 wuc1 = 2.527447264e-15 puc1 = -1.582749922e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.095525005e-01 lvth0 = -2.073743924e-07 wvth0 = -3.878494611e-07 pvth0 = 2.706763360e-13
+ k1 = -8.181497841e-01 lk1 = 7.650084241e-07 wk1 = 1.716588442e-06 pk1 = -9.864183589e-13
+ k2 = 5.198290321e-01 lk2 = -2.866642327e-07 wk2 = -7.017034236e-07 pk2 = 3.829158503e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.051200765e+00 ldsub = -1.751327196e-06 wdsub = -9.551422486e-06 pdsub = 2.622918174e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.104709678e-02 lvoff = -1.127513979e-07 wvoff = -2.894302384e-07 pvoff = 1.497864447e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -3.588867805e+00 lnfactor = 9.453451281e-07 wnfactor = 9.361741204e-06 pnfactor = -1.363937944e-12
+ eta0 = -3.024975615e+00 leta0 = 8.396222251e-07 weta0 = 4.589229492e-06 peta0 = -1.096229249e-12
+ etab = 2.418731793e-03 letab = -1.221856194e-09 wetab = -4.745851160e-09 petab = 1.972635199e-15
+ u0 = 1.566285551e-02 lu0 = -6.132845377e-09 wu0 = -5.834461978e-09 pu0 = 7.110373971e-15
+ ua = -1.685710765e-09 lua = -8.085154534e-16 wua = 2.109523131e-15 pua = 7.713518487e-22
+ ub = 4.199311452e-18 lub = -5.196496039e-25 wub = -4.902543649e-24 pub = 1.062239223e-30
+ uc = -4.240296082e-11 luc = 1.445267744e-18 wuc = -2.059901347e-17 puc = 1.627274566e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.843229381e+05 lvsat = -1.799723191e-02 wvsat = -2.139134616e-01 pvsat = 3.893139061e-8
+ a0 = 4.093929001e+00 la0 = -6.648828128e-07 wa0 = -4.255730168e-06 pa0 = 7.928346043e-13
+ ags = 2.162616775e+00 lags = -4.399870593e-07 wags = -1.537837347e-06 pags = 7.437548161e-13
+ a1 = 0.0
+ a2 = 1.825532881e+00 la2 = -3.873803105e-07 wa2 = -8.536367079e-07 pa2 = 3.898434891e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.456765088e-02 lketa = -5.987495946e-08 wketa = -1.129304222e-07 pketa = 8.086112170e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.841918725e+00 lpclm = -9.042380533e-07 wpclm = -7.047250150e-06 ppclm = 1.553058645e-12
+ pdiblc1 = 7.820230090e+00 lpdiblc1 = -1.715595191e-06 wpdiblc1 = -1.069214971e-05 ppdiblc1 = 2.482519326e-12
+ pdiblc2 = -3.245454199e-03 lpdiblc2 = 3.683721488e-09 wpdiblc2 = -7.128930104e-09 ppdiblc2 = 7.726965207e-16
+ pdiblcb = 3.656277649e-01 lpdiblcb = -1.474921849e-07 wpdiblcb = -2.571648646e-07 ppdiblcb = 7.245149502e-14
+ drout = 4.320364309e-01 ldrout = 2.165005493e-07 wdrout = 1.378934302e-06 pdrout = -5.942680310e-13
+ pscbe1 = 7.255521866e+08 lpscbe1 = 1.780650037e+01 wpscbe1 = 9.723681804e+01 ppscbe1 = -2.326621417e-5
+ pscbe2 = 8.037511926e-09 lpscbe2 = 4.383660503e-16 wpscbe2 = 1.901230561e-15 ppscbe2 = -6.780072136e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.310671459e+01 lbeta0 = -1.002000316e-06 wbeta0 = -5.942036353e-06 pbeta0 = 1.433320203e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.422210675e-09 lagidl = 5.926619789e-16 wagidl = 2.223773546e-15 pagidl = -8.302474840e-22
+ bgidl = 3.496250376e+09 lbgidl = -8.044895054e+02 wbgidl = -3.583967246e+03 pbgidl = 1.209148005e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.675370351e-01 lkt1 = -8.198862590e-08 wkt1 = -5.095546413e-07 pkt1 = 1.196485626e-13
+ kt2 = -1.576485041e-01 lkt2 = 2.935445787e-08 wkt2 = 1.885285464e-07 pkt2 = -5.071737710e-14
+ at = 2.573329861e+05 lat = -1.088408588e-01 wat = -3.362794043e-01 pat = 1.646494445e-7
+ ute = -1.551221188e+00 lute = 1.040785517e-06 wute = 2.596372332e-06 pute = -1.764778819e-12
+ ua1 = -1.127402449e-09 lua1 = 9.233371685e-16 wua1 = 7.662242818e-15 pua1 = -2.593628028e-21
+ ub1 = 3.127765906e-18 lub1 = -1.095234105e-24 wub1 = -1.009267066e-23 pub1 = 2.811068807e-30
+ uc1 = 4.591558542e-10 luc1 = -5.406471267e-17 wuc1 = -9.688805635e-16 puc1 = 1.264998632e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -2.666577256e+00 lvth0 = 2.786110244e-07 wvth0 = 2.591628106e-06 pvth0 = -4.724189824e-13
+ k1 = 7.210832963e+00 lk1 = -1.234922952e-06 wk1 = -1.059662811e-05 pk1 = 2.093962526e-12
+ k2 = -2.543023256e+00 lk2 = 4.766263424e-07 wk2 = 4.059876588e-06 pk2 = -8.081781119e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.332924860e+00 ldsub = 1.036889841e-06 wdsub = 8.300456742e-06 pdsub = -1.758173227e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.624848584e+00 lvoff = 2.895889502e-07 wvoff = 2.256706096e-06 pvoff = -4.910333948e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.754245750e+00 lnfactor = -3.545186200e-07 wnfactor = 1.302426625e-06 pnfactor = 6.011295715e-13
+ eta0 = -2.416206241e+00 leta0 = 7.436109908e-07 weta0 = 4.927827239e-06 peta0 = -1.260883156e-12
+ etab = -2.396507037e-01 letab = 6.062949270e-08 wetab = 4.052972418e-07 petab = -1.028047017e-13
+ u0 = -4.999103732e-02 lu0 = 1.022955128e-08 wu0 = 9.172234514e-08 pu0 = -1.734545220e-14
+ ua = -1.416655940e-08 lua = 2.327418522e-15 wua = 2.076223657e-14 pua = -3.946422049e-21
+ ub = 3.502293763e-18 lub = -3.782863280e-25 wub = -2.962470612e-24 pub = 6.414306201e-31
+ uc = -1.827144559e-10 luc = 3.744962740e-17 wuc = 2.956993542e-16 puc = -6.350041211e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.507911992e+04 lvsat = 3.686033815e-02 wvsat = 1.933373938e-01 pvsat = -6.250120029e-8
+ a0 = 1.895212042e+00 la0 = -1.496157623e-07 wa0 = -1.928112195e-06 pa0 = 2.536917781e-13
+ ags = -2.146985229e+00 lags = 6.313976225e-07 wags = 5.760002842e-06 pags = -1.070611699e-12
+ a1 = 0.0
+ a2 = -1.120302326e+00 la2 = 3.388013000e-07 wa2 = 3.023593805e-06 pa2 = -5.744789379e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.324608183e-01 lketa = 3.233410879e-08 wketa = 4.398592993e-07 pketa = -5.482642622e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.798236115e+00 lpclm = -1.898041755e-07 wpclm = -1.803371477e-06 ppclm = 3.218361356e-13
+ pdiblc1 = 4.213889025e-01 lpdiblc1 = 5.545010798e-08 wpdiblc1 = 6.807510406e-08 ppdiblc1 = -9.402242300e-14
+ pdiblc2 = 3.004518231e-04 lpdiblc2 = 3.038595145e-09 wpdiblc2 = 1.624230093e-08 ppdiblc2 = -5.152308776e-15
+ pdiblcb = -3.275013682e-01 lpdiblcb = 1.936198095e-08 wpdiblcb = 1.744541379e-07 ppdiblcb = -3.283060087e-14
+ drout = 2.603263332e+00 ldrout = -3.236432763e-07 wdrout = -3.253643984e-06 pdrout = 5.487766594e-13
+ pscbe1 = 8.003542628e+08 lpscbe1 = -6.584640191e-02 wpscbe1 = -6.006948682e-01 ppscbe1 = 1.116506077e-7
+ pscbe2 = 1.055147437e-08 lpscbe2 = -1.736837026e-16 wpscbe2 = -2.088146159e-15 ppscbe2 = 2.945019071e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.269033156e+00 lbeta0 = 1.187986454e-06 wbeta0 = 7.931037088e-06 pbeta0 = -2.014375967e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.481786397e-08 lagidl = -3.520507105e-15 wagidl = -2.458196446e-14 pagidl = 5.969449299e-21
+ bgidl = -2.186116388e+09 lbgidl = 5.922034331e+02 wbgidl = 5.402449000e+03 pbgidl = -1.004153170e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.505532930e-01 lkt1 = 6.135274321e-08 wkt1 = 3.979172103e-07 pkt1 = -1.040310612e-13
+ kt2 = -3.615905713e-02 lkt2 = 3.580634082e-10 wkt2 = -2.142069499e-08 pkt2 = -6.071401923e-16
+ at = -5.786981700e+05 lat = 9.732840140e-02 wat = 9.979898092e-01 pat = -1.650321786e-7
+ ute = 8.007161163e+00 lute = -1.330846717e-06 wute = -1.361103106e-05 pute = 2.256612971e-12
+ ua1 = 3.983878706e-09 lua1 = -3.187738951e-16 wua1 = -5.308142382e-15 pua1 = 5.405200295e-22
+ ub1 = -1.170777320e-18 lub1 = -7.331192822e-26 wub1 = 1.189694635e-24 pub1 = 1.243093183e-31
+ uc1 = 6.884804967e-10 luc1 = -1.165897090e-16 wuc1 = -1.211931399e-15 puc1 = 1.976920756e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.916867486e-01 lvth0 = -6.987487426e-08 wvth0 = -4.408631809e-07 pvth0 = 9.123017308e-14
+ k1 = -2.310853057e+00 lk1 = 5.348728284e-07 wk1 = 4.426260242e-06 pk1 = -6.983417319e-13
+ k2 = 1.379903914e+00 lk2 = -2.525281308e-07 wk2 = -2.062060224e-06 pk2 = 3.297062832e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.264155629e+00 ldsub = -1.118659509e-06 wdsub = -9.016591154e-06 pdsub = 1.460546466e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.742863937e+00 lvoff = -3.363677762e-07 wvoff = -2.747880785e-06 pvoff = 4.391691687e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -2.496859299e+01 lnfactor = 4.612455416e-06 wnfactor = 3.693621818e-05 pnfactor = -6.022123265e-12
+ eta0 = 9.214556518e+00 leta0 = -1.418198883e-06 weta0 = -1.181782735e-05 peta0 = 1.851631662e-12
+ etab = 1.098339872e+00 letab = -1.880628155e-07 wetab = -1.468827959e-06 petab = 2.455389493e-13
+ u0 = 1.452197892e-02 lu0 = -1.761483049e-09 wu0 = -1.397132905e-08 pu0 = 2.299831022e-15
+ ua = -2.554588734e-11 lua = -3.009716603e-16 wua = -2.584066058e-15 pua = 3.929552211e-22
+ ub = 8.793904358e-19 lub = 1.092327134e-25 wub = 1.255785448e-24 pub = -1.426166337e-31
+ uc = 9.799438381e-11 luc = -1.472572463e-17 wuc = -1.493786151e-16 puc = 1.922623004e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.025358830e+05 lvsat = -6.306616245e-02 wvsat = -5.859264435e-01 pvsat = 8.234056915e-8
+ a0 = 3.454250056e+00 la0 = -4.393941580e-07 wa0 = -3.649696643e-06 pa0 = 5.736826794e-13
+ ags = 1.249999265e+00 lags = 1.145400343e-13 wags = 9.594276591e-13 pags = -1.495459898e-19
+ a1 = 0.0
+ a2 = -1.061225533e-01 la2 = 1.502957057e-07 wa2 = 9.885717038e-07 pa2 = -1.962293799e-13
+ b0 = -4.760275983e-23 lb0 = 8.847924970e-30 wb0 = 6.215121049e-29 pb0 = -1.155204549e-35
+ b1 = 0.0
+ keta = -1.407787164e+00 lketa = 2.322050167e-07 wketa = 1.775984291e-06 pketa = -3.031719784e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.315397010e+00 lpclm = -2.859288711e-07 wpclm = -2.080333273e-06 ppclm = 3.733150245e-13
+ pdiblc1 = 7.394020791e+00 lpdiblc1 = -1.240552981e-06 wpdiblc1 = -9.151894161e-06 ppdiblc1 = 1.619693264e-12
+ pdiblc2 = 1.492542833e-01 lpdiblc2 = -2.464745351e-08 wpdiblc2 = -1.846108024e-07 ppdiblc2 = 3.218025754e-14
+ pdiblcb = -3.603082878e+00 lpdiblcb = 6.281943163e-07 wpdiblcb = 4.410499324e-06 ppdiblcb = -8.201843196e-13
+ drout = -6.266896325e+00 ldrout = 1.325053299e-06 wdrout = 9.006513105e-06 pdrout = -1.730018739e-12
+ pscbe1 = 8.084381355e+08 lpscbe1 = -1.568395831e+00 wpscbe1 = -1.101701538e+01 ppscbe1 = 2.047732102e-6
+ pscbe2 = 4.474533569e-08 lpscbe2 = -6.529296706e-15 wpscbe2 = -4.636797355e-14 ppscbe2 = 8.524793424e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.627803013e+01 lbeta0 = -2.902825813e-06 wbeta0 = -2.329707509e-05 pbeta0 = 3.789993244e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.202834507e-08 lagidl = 1.469397768e-15 wagidl = 1.785590799e-14 pagidl = -1.918478053e-21
+ bgidl = 9.999993372e+08 lbgidl = 1.033171067e-04 wbgidl = 8.654204636e-04 pbgidl = -1.348930874e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.233304002e-01 lkt1 = -1.196630188e-07 wkt1 = -1.002339588e-06 pkt1 = 1.562346700e-13
+ kt2 = 6.400896291e-02 lkt2 = -1.826016648e-08 wkt2 = -1.529535689e-07 pkt2 = 2.384087508e-14
+ at = -4.931973912e+05 lat = 8.143637166e-02 wat = 6.821396978e-01 pat = -1.063251184e-7
+ ute = 6.697734947e+00 lute = -1.087463666e-06 wute = -9.108978634e-06 pute = 1.419816486e-12
+ ua1 = 1.074914996e-08 lua1 = -1.576234863e-15 wua1 = -1.347216501e-14 pua1 = 2.057966915e-21
+ ub1 = -8.960991806e-18 lub1 = 1.374655238e-24 wub1 = 1.151459612e-23 pub1 = -1.794780121e-30
+ uc1 = 6.514783155e-10 luc1 = -1.097121136e-16 wuc1 = -9.189872634e-16 puc1 = 1.432425492e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.071200549e+00 lvth0 = 1.888858026e-07 wvth0 = -3.152484594e-08 pvth0 = 6.301460472e-13
+ k1 = 1.059737551e+00 lk1 = -1.223758322e-05 wk1 = -7.367258537e-07 pk1 = 1.472631731e-11
+ k2 = -8.856083998e-02 lk2 = 2.199954043e-06 wk2 = 1.250090640e-07 pk2 = -2.498789929e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.106833681e-04 lcit = -2.012546757e-09 wcit = -1.314544205e-10 pcit = 2.627625322e-15
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.701450401e-02 lvoff = -5.400281550e-06 wvoff = -3.685321472e-07 pvoff = 7.366541181e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -4.858103329e+00 lnfactor = 1.399362067e-04 wnfactor = 8.165812788e-06 pnfactor = -1.632253703e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.610096683e-02 lu0 = -5.303340414e-07 wu0 = -2.897754111e-08 pu0 = 5.792283021e-13
+ ua = 1.386374813e-09 lua = -4.084291533e-14 wua = -2.591034058e-15 pua = 5.179184294e-20
+ ub = 4.464896017e-18 lub = -6.876760766e-23 wub = -3.444946661e-24 pub = 6.886059097e-29
+ uc = -1.553851903e-10 luc = 1.671235065e-15 wuc = 4.808819537e-17 puc = -9.612286857e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.944361679e+05 lvsat = -1.667323953e+01 wvsat = -1.089049396e+00 pvsat = 2.176886680e-5
+ a0 = 3.305086701e+00 la0 = -3.918623474e-05 wa0 = -2.111261173e-06 pa0 = 4.220172512e-11
+ ags = 4.378176839e+00 lags = -8.449812738e-05 wags = -4.982204831e-06 pags = 9.958864468e-11
+ a1 = 0.0
+ a2 = -9.690507613e-01 la2 = 3.536132569e-05 wa2 = 2.309711593e-06 pa2 = -4.616852477e-11
+ b0 = 1.070067587e-06 lb0 = -2.138944189e-11 wb0 = -1.397103783e-12 pb0 = 2.792652590e-17
+ b1 = -2.411944620e-08 lb1 = 4.821204746e-13 wb1 = 3.149087959e-14 pb1 = -6.294670983e-19
+ keta = -6.067220295e-01 lketa = 1.209030459e-05 wketa = 7.417874372e-07 pketa = -1.482749265e-11
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.097533665e-01 lpclm = -7.371783048e-06 wpclm = -6.133801217e-07 ppclm = 1.226077551e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.002496346e-02 lpdiblc2 = 2.067700979e-07 wpdiblc2 = 1.345297292e-08 ppdiblc2 = -2.689097267e-13
+ pdiblcb = 2.362311511e+00 lpdiblcb = -5.032060181e-05 wpdiblcb = -3.036179439e-06 ppdiblcb = 6.068979610e-11
+ drout = 0.56
+ pscbe1 = 6.864776709e+08 lpscbe1 = 2.268208620e+03 wpscbe1 = 1.323383224e+02 ppscbe1 = -2.645293522e-3
+ pscbe2 = 3.058498191e-09 lpscbe2 = 4.731294787e-14 wpscbe2 = 9.511793143e-15 ppscbe2 = -1.901299966e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.140618095e-09 lalpha0 = -2.080077982e-14 walpha0 = -1.358653878e-15 palpha0 = 2.715795575e-20
+ alpha1 = 1.140618095e-09 lalpha1 = -2.080077982e-14 walpha1 = -1.358653878e-15 palpha1 = 2.715795575e-20
+ beta0 = -2.787860768e+02 lbeta0 = 5.698120552e-03 wbeta0 = 3.668365471e-04 pbeta0 = -7.332648052e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.818464735e-08 lagidl = 3.723875525e-13 wagidl = 2.383521239e-14 pagidl = -4.764389620e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.625313682e-02 legidl = 1.962312938e-05 pegidl = 7.105427358e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.391529389e-01 lkt1 = 3.965420793e-06 wkt1 = 2.349112556e-07 pkt1 = -4.695610549e-12
+ kt2 = 1.798475998e-01 lkt2 = -4.641536982e-06 wkt2 = -2.796789008e-07 pkt2 = 5.590465191e-12
+ at = -7.387347856e+05 lat = 1.476647359e+01 wat = 9.645083882e-01 pat = -1.927943279e-5
+ ute = -2.946327405e+00 lute = 5.624990520e-05 wute = 3.351934983e-06 pute = -6.700139263e-11
+ ua1 = 6.923187214e-09 lua1 = -1.019524901e-13 wua1 = -5.555535708e-15 pua1 = 1.110488811e-19
+ ub1 = -6.624446708e-18 lub1 = 1.181053943e-22 wub1 = 6.139756876e-24 pub1 = -1.227268020e-28
+ uc1 = 5.276253915e-09 luc1 = -1.056414815e-13 wuc1 = -6.190964541e-15 puc1 = 1.237503854e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.061751
+ k1 = 0.44751769
+ k2 = 0.02149811
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.23314992
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1426029
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0095695
+ ua = -6.5690804e-10
+ ub = 1.02460111e-18
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.344684
+ ags = 0.150918
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-01 pvsat = -1.862645149e-21
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595752e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 ppdiblc2 = -6.938893904e-30
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+3
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 wpscbe2 = -1.323488980e-29
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17 wuc1 = -2.584939414e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569066e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16 wua = 1.654361225e-30
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077653e-03 lketa = -3.715224604e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = 2.220446049e-22 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048849e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807946e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-02 wat = -2.328306437e-16
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123885e-18 lub1 = 2.335179770e-24 wub1 = 6.162975822e-39
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-08 pk2 = -1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = -1.058181320e-22 peta0 = -3.191891196e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = -6.817463261e-22 petab = 7.580741590e-28
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-09 wu0 = 2.775557562e-23
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16 pagidl = 8.271806126e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = 6.661338148e-22 pute = -8.881784197e-28
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24 wub1 = 6.162975822e-39 pub1 = 6.162975822e-45
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 wuc1 = 1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.68 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.059631612e+00 lvth0 = 2.586054434e-8
+ k1 = 5.163379589e-01 lk1 = -1.485963682e-10
+ k2 = -3.690874683e-03 lk2 = -1.907482336e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.279561642e+00 ldsub = -4.971871951e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.986924020e-01 lvoff = -1.955441768e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.816966235e+00 lnfactor = 7.632892377e-7
+ eta0 = -4.398980000e-02 leta0 = 2.610515935e-7
+ etab = -1.632772774e+00 letab = 7.979080824e-7
+ u0 = 8.012298384e-03 lu0 = 8.686250060e-10
+ ua = -7.759682813e-10 lua = 1.274097302e-16
+ ub = 6.727035311e-19 lub = 1.823100696e-25
+ uc = -9.895092236e-11 luc = 3.384048354e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.003651958e+04 lvsat = -2.626952517e-03 wvsat = -1.164153218e-16
+ a0 = 1.678264962e+00 la0 = -4.701829257e-7
+ ags = -3.625107542e-01 lags = 7.883081324e-07 pags = -8.881784197e-28
+ a1 = 0.0
+ a2 = 1.009669841e+00 la2 = -9.572104471e-9
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.793248020e-03 lketa = -2.322682382e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.567025060e+00 lpclm = -7.524585059e-7
+ pdiblc1 = 6.637643939e-02 lpdiblc1 = -2.707173962e-8
+ pdiblc2 = 8.111861681e-04 lpdiblc2 = -3.769435660e-10
+ pdiblcb = -3.034907083e-02 lpdiblcb = 5.289535676e-9
+ drout = 1.0
+ pscbe1 = 7.729094317e+08 lpscbe1 = 1.324376613e+1
+ pscbe2 = 9.028731239e-09 lpscbe2 = 1.463768495e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.609000049e+00 lbeta0 = 1.047440030e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.165212580e-10 lagidl = -3.050311102e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.213729371e-01 lkt1 = -5.704969315e-8
+ kt2 = -6.409955753e-02 lkt2 = 1.536741214e-8
+ at = 8.783879526e+04 lat = -2.578681467e-2
+ ute = -1.878857286e+00 lute = 8.214518228e-7
+ ua1 = -3.360596897e-09 lua1 = 2.897579860e-15 wua1 = -1.654361225e-30 pua1 = -3.308722450e-36
+ ub1 = 4.154167712e-18 lub1 = -3.223006351e-24 wub1 = -3.081487911e-39 pub1 = -3.081487911e-45
+ uc1 = 3.233299061e-10 luc1 = -2.535572683e-16 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.69 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.006613565e+00 lvth0 = -5.838818845e-11
+ k1 = 4.966170030e-01 lk1 = 9.492387336e-9
+ k2 = -1.761857806e-02 lk2 = 6.618088114e-09 wk2 = -1.387778781e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.644100980e-01 ldsub = 2.576142694e-07 pdsub = 2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.427270611e-01 lvoff = 1.972806098e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.581462661e+00 lnfactor = -9.932013026e-8
+ eta0 = 0.49
+ etab = -1.216203250e-03 letab = 2.890215328e-10
+ u0 = 1.119413334e-02 lu0 = -6.868786489e-10
+ ua = -6.998804391e-11 lua = -2.177228284e-16
+ ub = 4.443627388e-19 lub = 2.939390328e-25
+ uc = -5.818012563e-11 luc = 1.390886414e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.048266764e+04 lvsat = 1.182103908e-2
+ a0 = 8.343866772e-01 la0 = -5.763614858e-8
+ ags = 9.847587520e-01 lags = 1.296684889e-7
+ a1 = 0.0
+ a2 = 1.171716763e+00 la2 = -8.879198318e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.192784488e-02 lketa = 2.058066866e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.557003024e-01 lpclm = 2.852782422e-07 wpclm = -1.110223025e-22 ppclm = 8.326672685e-29
+ pdiblc1 = -3.690848156e-01 lpdiblc1 = 1.858122041e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = 1.249000903e-28
+ pdiblc2 = -8.705633412e-03 lpdiblc2 = 4.275544022e-09 wpdiblc2 = -1.626303259e-24 ppdiblc2 = 8.673617380e-31
+ pdiblcb = 1.686604462e-01 lpdiblcb = -9.200024691e-08 wpdiblcb = 1.110223025e-22 ppdiblcb = 1.110223025e-28
+ drout = 1.488187677e+00 ldrout = -2.386603096e-07 wdrout = 3.552713679e-21
+ pscbe1 = 8.000276611e+08 lpscbe1 = -1.352270444e-02 wpscbe1 = -1.907348633e-12
+ pscbe2 = 9.493699522e-09 lpscbe2 = -8.093219498e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.555599215e+00 lbeta0 = 9.580609553e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.810185489e-10 lagidl = -4.323990079e-17
+ bgidl = 7.512236789e+08 lbgidl = 1.216192801e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.578143445e-01 lkt1 = 9.652417683e-9
+ kt2 = -1.325100891e-02 lkt2 = -9.490917822e-9
+ at = -2.296195638e+02 lat = 1.726719129e-2
+ ute = 4.373883268e-01 lute = -3.108911698e-07 pute = -2.220446049e-28
+ ua1 = 4.741250820e-09 lua1 = -1.063170433e-15
+ ub1 = -4.602396930e-18 lub1 = 1.057815405e-24
+ uc1 = -2.829276611e-10 luc1 = 4.282386859e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.70 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.506813703e-01 lvth0 = -2.045149115e-07 wvth0 = -7.320212644e-07 pvth0 = 1.748579194e-13
+ k1 = -3.489492597e+00 lk1 = 9.616543876e-07 wk1 = 3.546109364e-06 pk1 = -8.470591438e-13
+ k2 = 1.907088917e+00 lk2 = -4.531367913e-07 wk2 = -1.816732860e-06 pk2 = 4.339629783e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.480511613e+01 ldsub = -3.342043460e-06 wdsub = -1.683114040e-05 pdsub = 4.020454508e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.924900471e-01 lvoff = -1.497615045e-07 wvoff = -4.175463558e-07 pvoff = 9.973929801e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -4.333466577e+00 lnfactor = 1.791319017e-06 wnfactor = 9.300100178e-06 pnfactor = -2.221514930e-12
+ eta0 = 6.192648726e+00 leta0 = -1.362191701e-06 weta0 = -6.415747845e-06 peta0 = 1.532529688e-12
+ etab = 5.997079623e-01 letab = -1.432537339e-07 wetab = -6.990400796e-07 petab = 1.669797038e-13
+ u0 = 2.773946023e-02 lu0 = -4.639060883e-09 wu0 = -1.119037451e-08 pu0 = 2.673044758e-15
+ ua = 3.242098858e-09 lua = -1.008881027e-15 wua = -2.291349287e-15 pua = 5.473346041e-22
+ ub = 4.221177318e-18 lub = -6.082286659e-25 wub = -3.848325001e-24 pub = 9.192493931e-31
+ uc = 1.720747195e-10 luc = -4.109211072e-17 wuc = -1.727419421e-16 puc = 4.126286772e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.131855634e+05 lvsat = -1.775319016e-01 wvsat = -9.193142310e-01 pvsat = 2.195965904e-7
+ a0 = 5.590577153e+00 la0 = -1.193747368e-06 wa0 = -6.732004685e-06 pa0 = 1.608073959e-12
+ ags = 2.197290171e+00 lags = -1.599688912e-7
+ a1 = 0.0
+ a2 = -4.779319936e-01 la2 = 3.052596153e-07 wa2 = 2.137669664e-06 pa2 = -5.106251527e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.672537229e-02 lketa = 7.981452239e-09 wketa = 8.840165087e-08 pketa = -2.111650234e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.339806916e-01 lpclm = 2.323160788e-07 wpclm = 1.006957741e-06 ppclm = -2.405319957e-13
+ pdiblc1 = 7.463804736e-01 lpdiblc1 = -8.063898952e-08 wpdiblc1 = -3.639711791e-07 ppdiblc1 = 8.694179555e-14
+ pdiblc2 = 5.420951848e-02 lpdiblc2 = -1.075299831e-08 wpdiblc2 = -5.456616419e-08 ppdiblc2 = 1.303421964e-14
+ pdiblcb = 1.638952311e+00 lpdiblcb = -4.432088647e-07 wpdiblcb = -2.395690246e-06 ppdiblcb = 5.722585289e-13
+ drout = -2.702161725e+00 ldrout = 7.622884521e-07 wdrout = 3.718353858e-06 pdrout = -8.882031860e-13
+ pscbe1 = 7.999012102e+08 lpscbe1 = 1.668263473e-2
+ pscbe2 = -4.273794744e-08 lpscbe2 = 1.239564132e-14 wpscbe2 = 6.751190807e-14 ppscbe2 = -1.612656948e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.672541998e+01 lbeta0 = -4.244418991e-06 wbeta0 = -2.155412933e-05 pbeta0 = 5.148634872e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.221889522e-08 lagidl = 7.720014502e-15 wagidl = 3.732104681e-14 pagidl = -8.914878451e-21
+ bgidl = 1.888486861e+09 lbgidl = -1.500387762e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.318186390e-01 lkt1 = -4.433117647e-08 wkt1 = -1.573449734e-07 pkt1 = 3.758499379e-14
+ kt2 = 1.509835437e-01 lkt2 = -4.872162540e-08 wkt2 = -2.658081083e-07 pkt2 = 6.349358284e-14
+ at = 6.155641632e+05 lat = -1.298274696e-01 wat = -5.748336360e-01 pat = 1.373105106e-7
+ ute = -1.647000087e+00 lute = 1.870066905e-07 wute = -8.208162777e-07 pute = 1.960683843e-13
+ ua1 = -4.787079780e-09 lua1 = 1.212861897e-15 wua1 = 6.187853319e-15 pua1 = -1.478092522e-21
+ ub1 = 9.994511496e-18 lub1 = -2.428948111e-24 wub1 = -1.337773188e-23 pub1 = 3.195538813e-30
+ uc1 = 1.189237198e-10 luc1 = -5.316637077e-17 wuc1 = -4.520521085e-16 puc1 = 1.079816871e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.71 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -2.651426023e+00 lvth0 = 2.397101539e-07 wvth0 = 1.987253330e-06 pvth0 = -3.129708506e-13
+ k1 = 7.999139645e+00 lk1 = -1.076928754e-06 wk1 = -9.034693050e-06 pk1 = 1.406061874e-12
+ k2 = -3.794094283e+00 lk2 = 5.609252328e-07 wk2 = 4.693225651e-06 pk2 = -7.323563243e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -3.515572503e+01 ldsub = 5.607737399e-06 wdsub = 4.636773827e-05 pdsub = -7.321585318e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.551677196e+00 lvoff = 1.965244971e-07 wvoff = 1.553544598e-06 pvoff = -2.565867069e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.487234672e+01 lnfactor = -3.456834931e-06 wnfactor = -2.813720920e-05 pnfactor = 4.513319736e-12
+ eta0 = -1.077748539e+01 leta0 = 1.654916441e-06 weta0 = 1.428422239e-05 peta0 = -2.160695313e-12
+ etab = -7.488466977e-01 letab = 9.298088860e-08 wetab = 9.428994643e-07 petab = -1.213978937e-13
+ u0 = -1.317212355e-02 lu0 = 2.498164860e-09 wu0 = 2.218670040e-08 pu0 = -3.261659001e-15
+ ua = -4.463787585e-09 lua = 3.218488872e-16 wua = 3.210599943e-15 pua = -4.202129878e-22
+ ub = -5.868961389e-18 lub = 1.205995551e-24 wub = 1.006658205e-23 pub = -1.574574323e-30
+ uc = 3.546895544e-10 luc = -7.917143810e-17 wuc = -4.845254772e-16 puc = 1.033679714e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.832960690e+06 lvsat = 2.964353161e-01 wvsat = 2.463349263e+00 pvsat = -3.870324703e-7
+ a0 = -1.425669903e+00 la0 = -9.811064619e-09 wa0 = 2.721634213e-06 pa0 = 1.280954181e-14
+ ags = 1.25
+ a1 = 0.0
+ a2 = 1.158116137e+01 la2 = -1.905433840e-06 wa2 = -1.427060330e-05 pa2 = 2.487776341e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.159744099e+00 lketa = -4.050489423e-07 wketa = -2.881863012e-06 pketa = 5.288408101e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.614603622e+00 lpclm = 4.937325259e-07 wpclm = 3.050762012e-06 ppclm = -6.446280479e-13
+ pdiblc1 = -1.033719298e+01 lpdiblc1 = 1.971346950e-06 wpdiblc1 = 1.399836863e-05 ppdiblc1 = -2.573833947e-12
+ pdiblc2 = -3.167657868e-01 lpdiblc2 = 5.711768644e-08 wpdiblc2 = 4.238352535e-07 ppdiblc2 = -7.457410800e-14
+ pdiblcb = -9.803990370e+00 lpdiblcb = 1.639073430e-06 wpdiblcb = 1.250654056e-05 ppdiblcb = -2.140010330e-12
+ drout = 2.389245913e+01 ldrout = -4.104114793e-06 wdrout = -3.037020488e-05 pdrout = 5.358422564e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 1.033768946e-07 lpscbe2 = -1.351486566e-14 wpscbe2 = -1.229186268e-13 ppscbe2 = 1.764530594e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -4.282785357e+01 lbeta0 = 8.256165896e-06 wbeta0 = 6.692908699e-05 pbeta0 = -1.077943183e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.698085916e-08 lagidl = -2.506276518e-15 wagidl = -3.307536725e-14 pagidl = 3.272249760e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.800812639e+00 lkt1 = 2.242479564e-07 wkt1 = 1.640426096e-06 pkt1 = -2.927830653e-13
+ kt2 = -2.441216247e+00 lkt2 = 4.281857850e-07 wkt2 = 3.117923581e-06 pkt2 = -5.590487809e-13
+ at = -1.404574883e+06 lat = 2.325861534e-01 wat = 1.872054201e+00 pat = -3.036695988e-7
+ ute = 9.959223438e+00 lute = -1.951416271e-06 wute = -1.336724976e-05 pute = 2.547812014e-12
+ ua1 = 2.614271089e-08 lua1 = -4.413960513e-15 wua1 = -3.357033681e-14 pua1 = 5.762963953e-21
+ ub1 = -4.076849220e-17 lub1 = 6.761851236e-24 wub1 = 5.304316841e-23 pub1 = -8.828421735e-30
+ uc1 = 3.757067888e-10 luc1 = -1.062468534e-16 wuc1 = -5.589338911e-16 puc1 = 1.387182292e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.72 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.098246063e+00 lvth0 = 7.294950629e-7
+ k1 = 4.276922968e-01 lk1 = 3.962872071e-07 wk1 = 8.881784197e-22
+ k2 = 1.868581804e-02 lk2 = 5.621453833e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.092832443e-06 lcit = 2.417220556e-10 wcit = -1.694065895e-27 pcit = 1.761828530e-31
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.791532993e-01 lvoff = 9.195555675e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.147437737e+00 lnfactor = -9.664292472e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.124081396e-02 lu0 = -3.340767752e-8
+ ua = -8.365019490e-10 lua = 3.589879299e-15
+ ub = 1.509438192e-18 lub = -9.691345396e-24
+ uc = -1.141297958e-10 luc = 8.465863493e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.012865143e+04 lvsat = 2.002511953e+0
+ a0 = 1.493812400e+00 la0 = -2.980908204e-6
+ ags = 1.038882350e-01 lags = 9.400718588e-7
+ a1 = 0.0
+ a2 = 1.012476349e+00 la2 = -4.247162113e-06 wa2 = -1.776356839e-21
+ b0 = -1.285231938e-07 lb0 = 2.569033412e-12
+ b1 = 2.896927536e-09 lb1 = -5.790630792e-14
+ keta = 2.966561342e-02 lketa = -6.303652749e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.647222096e-02 lpclm = 3.146871810e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.516490733e-03 lpdiblc2 = -2.393052950e-8
+ pdiblcb = -2.424603954e-01 lpdiblcb = 1.745845204e-6
+ drout = 0.56
+ pscbe1 = 8.000121807e+08 lpscbe1 = -1.217936194e+0
+ pscbe2 = 1.121877068e-08 lpscbe2 = -1.158016781e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.498608750e-11 lalpha0 = 2.498330655e-15
+ alpha1 = -2.498608750e-11 lalpha1 = 2.498330655e-15
+ beta0 = 3.592705243e+01 lbeta0 = -5.926392753e-04 pbeta0 = 9.094947018e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.263844868e-09 lagidl = -3.635470011e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.625313682e-02 legidl = 1.962312938e-05 pegidl = 1.065814104e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.376199758e-01 lkt1 = -6.299540746e-8
+ kt2 = -6.009202116e-02 lkt2 = 1.545849088e-7
+ at = 8.872762352e+04 lat = -1.773564932e+0
+ ute = -7.066532693e-02 lute = -1.231330245e-6
+ ua1 = 2.157031712e-09 lua1 = -6.682427407e-15
+ ub1 = -1.357081407e-18 lub1 = 1.281671407e-23
+ uc1 = -3.504300659e-11 luc1 = 5.253421821e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.73 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.061751
+ k1 = 0.44751769
+ k2 = 0.02149811
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.23314992
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1426029
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0095695
+ ua = -6.5690804e-10
+ ub = 1.02460111e-18
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.344684
+ ags = 0.150918
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.74 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-1
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595752e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-07 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 wpdiblc2 = 8.673617380e-25
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+03 wpscbe1 = -1.907348633e-12 ppscbe1 = -7.629394531e-18
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 wpscbe2 = 1.323488980e-29 ppscbe2 = -5.293955920e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23 pub1 = 1.232595164e-44
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.75 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569066e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077653e-03 lketa = -3.715224604e-08 wketa = 6.938893904e-24 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = 2.220446049e-22 ppclm = 1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048848e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807947e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123885e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.76 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = -1.734723476e-22 peta0 = -2.255140519e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = 7.424616477e-22 petab = -1.058181320e-27
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-9
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16 pagidl = -8.271806126e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = 4.440892099e-22 pute = 1.554312234e-27
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15 pua1 = -6.617444900e-36
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 wuc1 = 1.033975766e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.77 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.059631612e+00 lvth0 = 2.586054434e-8
+ k1 = 5.163379589e-01 lk1 = -1.485963682e-10
+ k2 = -3.690874683e-03 lk2 = -1.907482336e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.279561642e+00 ldsub = -4.971871951e-07 pdsub = -8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.986924020e-01 lvoff = -1.955441768e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.816966235e+00 lnfactor = 7.632892377e-7
+ eta0 = -4.398980000e-02 leta0 = 2.610515935e-7
+ etab = -1.632772774e+00 letab = 7.979080824e-7
+ u0 = 8.012298384e-03 lu0 = 8.686250060e-10
+ ua = -7.759682813e-10 lua = 1.274097302e-16
+ ub = 6.727035311e-19 lub = 1.823100696e-25
+ uc = -9.895092236e-11 luc = 3.384048354e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.003651958e+04 lvsat = -2.626952517e-3
+ a0 = 1.678264962e+00 la0 = -4.701829257e-7
+ ags = -3.625107542e-01 lags = 7.883081324e-07 pags = -8.881784197e-28
+ a1 = 0.0
+ a2 = 1.009669841e+00 la2 = -9.572104471e-9
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.793248020e-03 lketa = -2.322682382e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.567025060e+00 lpclm = -7.524585059e-7
+ pdiblc1 = 6.637643939e-02 lpdiblc1 = -2.707173962e-8
+ pdiblc2 = 8.111861681e-04 lpdiblc2 = -3.769435660e-10
+ pdiblcb = -3.034907083e-02 lpdiblcb = 5.289535676e-9
+ drout = 1.0
+ pscbe1 = 7.729094317e+08 lpscbe1 = 1.324376613e+1
+ pscbe2 = 9.028731239e-09 lpscbe2 = 1.463768495e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.609000049e+00 lbeta0 = 1.047440030e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.165212580e-10 lagidl = -3.050311102e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.213729371e-01 lkt1 = -5.704969315e-8
+ kt2 = -6.409955753e-02 lkt2 = 1.536741214e-8
+ at = 8.783879526e+04 lat = -2.578681467e-2
+ ute = -1.878857286e+00 lute = 8.214518228e-7
+ ua1 = -3.360596897e-09 lua1 = 2.897579860e-15 wua1 = 3.308722450e-30 pua1 = 1.654361225e-36
+ ub1 = 4.154167712e-18 lub1 = -3.223006351e-24
+ uc1 = 3.233299061e-10 luc1 = -2.535572683e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.78 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.006613565e+00 lvth0 = -5.838818845e-11
+ k1 = 4.966170030e-01 lk1 = 9.492387336e-9
+ k2 = -1.761857806e-02 lk2 = 6.618088114e-09 wk2 = -1.387778781e-23 pk2 = -3.469446952e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.644100980e-01 ldsub = 2.576142694e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.427270611e-01 lvoff = 1.972806098e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.581462661e+00 lnfactor = -9.932013026e-8
+ eta0 = 0.49
+ etab = -1.216203250e-03 letab = 2.890215328e-10
+ u0 = 1.119413334e-02 lu0 = -6.868786489e-10
+ ua = -6.998804391e-11 lua = -2.177228284e-16
+ ub = 4.443627388e-19 lub = 2.939390328e-25
+ uc = -5.818012563e-11 luc = 1.390886414e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.048266764e+04 lvsat = 1.182103908e-2
+ a0 = 8.343866772e-01 la0 = -5.763614858e-08 wa0 = -1.776356839e-21
+ ags = 9.847587520e-01 lags = 1.296684889e-7
+ a1 = 0.0
+ a2 = 1.171716763e+00 la2 = -8.879198318e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.192784488e-02 lketa = 2.058066866e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.557003024e-01 lpclm = 2.852782422e-07 wpclm = 3.330669074e-22 ppclm = 5.551115123e-29
+ pdiblc1 = -3.690848156e-01 lpdiblc1 = 1.858122041e-07 wpdiblc1 = 1.387778781e-22 ppdiblc1 = 9.020562075e-29
+ pdiblc2 = -8.705633412e-03 lpdiblc2 = 4.275544022e-09 wpdiblc2 = 2.059984128e-24 ppdiblc2 = -8.944667923e-31
+ pdiblcb = 1.686604462e-01 lpdiblcb = -9.200024691e-8
+ drout = 1.488187677e+00 ldrout = -2.386603096e-7
+ pscbe1 = 8.000276611e+08 lpscbe1 = -1.352270444e-2
+ pscbe2 = 9.493699522e-09 lpscbe2 = -8.093219498e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.555599215e+00 lbeta0 = 9.580609553e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.810185489e-10 lagidl = -4.323990079e-17
+ bgidl = 7.512236789e+08 lbgidl = 1.216192801e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.578143445e-01 lkt1 = 9.652417683e-9
+ kt2 = -1.325100891e-02 lkt2 = -9.490917822e-9
+ at = -2.296195638e+02 lat = 1.726719129e-2
+ ute = 4.373883268e-01 lute = -3.108911698e-07 wute = -4.440892099e-22 pute = 1.110223025e-28
+ ua1 = 4.741250820e-09 lua1 = -1.063170433e-15
+ ub1 = -4.602396930e-18 lub1 = 1.057815405e-24
+ uc1 = -2.829276611e-10 luc1 = 4.282386859e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.79 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.786905057e-01 lvth0 = -5.450236936e-8
+ k1 = -4.472461707e-01 lk1 = 2.349529836e-7
+ k2 = 3.484937124e-01 lk2 = -8.083515471e-08 wk2 = -1.665334537e-22 pk2 = -3.469446952e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.654947035e-01 ldsub = 1.071489094e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.427241235e-02 lvoff = -6.419405813e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.645192181e+00 lnfactor = -1.145432006e-7
+ eta0 = 6.885077223e-01 leta0 = -4.741753964e-8
+ etab = -6.25e-6
+ u0 = 1.813911423e-02 lu0 = -2.345826234e-9
+ ua = 1.276324974e-09 lua = -5.393166190e-16
+ ub = 9.196567555e-19 lub = 1.804055510e-25
+ uc = 2.387749767e-11 luc = -5.692240336e-18 wuc = 1.090521315e-32 puc = -1.918509721e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.449572143e+04 lvsat = 1.086244092e-2
+ a0 = -1.848840900e-01 la0 = 1.858370596e-7
+ ags = 2.197290171e+00 lags = -1.599688912e-7
+ a1 = 0.0
+ a2 = 1.355998444e+00 la2 = -1.328113483e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.115381286e-03 lketa = -1.013462857e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.298994868e-01 lpclm = 2.596102059e-8
+ pdiblc1 = 4.341255753e-01 lpdiblc1 = -6.050661960e-9
+ pdiblc2 = 7.396602975e-03 lpdiblc2 = 4.292028164e-10
+ pdiblcb = -4.163368351e-01 lpdiblcb = 4.773805368e-08 wpdiblcb = 8.881784197e-22
+ drout = 4.878551563e-01 ldrout = 2.891195681e-10
+ pscbe1 = 7.999012102e+08 lpscbe1 = 1.668263473e-2
+ pscbe2 = 1.518126485e-08 lpscbe2 = -1.439520925e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.233894147e+00 lbeta0 = 1.726517851e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.007565774e-10 lagidl = 7.184172364e-17
+ bgidl = 1.888486861e+09 lbgidl = -1.500387762e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.668066312e-01 lkt1 = -1.208659480e-8
+ kt2 = -7.705617102e-02 lkt2 = 5.750221250e-9
+ at = 1.224080320e+05 lat = -1.202726455e-2
+ ute = -2.351187446e+00 lute = 3.552159249e-7
+ ua1 = 5.215479907e-10 lua1 = -5.521001849e-17
+ ub1 = -1.482392574e-18 lub1 = 3.125399646e-25 wub1 = -7.703719778e-40
+ uc1 = -2.688967816e-10 luc1 = 3.947231239e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.80 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.465379578e-01 lvth0 = -2.879127084e-08 wvth0 = -1.706293730e-12 pvth0 = 3.171488174e-19
+ k1 = 2.481761779e-01 lk1 = 1.293473497e-07 wk1 = 4.892214349e-13 pk1 = -9.093158759e-20
+ k2 = 2.322757765e-01 lk2 = -6.737133359e-08 wk2 = 1.290675229e-13 pk2 = -2.398978061e-20
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.623670784e+00 ldsub = -6.735316886e-07 wdsub = -6.354215856e-13 pdsub = 1.181058096e-19
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.188749411e-01 lvoff = -2.360392105e-08 wvoff = 9.680344952e-13 pvoff = -1.799285716e-19
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.331236489e-01 lnfactor = 4.151920104e-07 wnfactor = 2.757657569e-13 pnfactor = -5.125657765e-20
+ eta0 = 1.477115255e+00 leta0 = -1.987695053e-07 weta0 = -9.719470487e-12 peta0 = 1.806557979e-18
+ etab = 6.007622203e-02 letab = -1.116752908e-08 wetab = 1.112744818e-12 petab = -2.068258792e-19
+ u0 = 5.862077829e-03 lu0 = -3.000458201e-10 wu0 = 1.652537224e-14 pu0 = -3.071570935e-21
+ ua = -1.709377372e-09 lua = -3.865667163e-17 wua = -1.198109707e-21 pua = 2.226926513e-28
+ ub = 2.767251528e-18 lub = -1.448456153e-25 wub = 2.228047492e-29 pub = -4.141271871e-36
+ uc = -6.099048795e-11 luc = 9.509139135e-18 wuc = 3.251912996e-22 puc = -6.044330686e-29
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.803741985e+05 lvsat = -3.560417888e-02 wvsat = -3.762949593e-07 pvsat = 6.994194398e-14
+ a0 = 9.092405073e-01 la0 = 1.180180203e-09 wa0 = 1.127111264e-11 pa0 = -2.094961706e-18
+ ags = 1.25
+ a1 = 0.0
+ a2 = -6.617445391e-01 la2 = 2.288565339e-07 wa2 = -2.834559893e-12 pa2 = 5.268596475e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.126349108e-01 lketa = 4.864885374e-08 wketa = -3.646202202e-12 pketa = 6.777196032e-19
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.002677566e+00 lpclm = -5.930076705e-08 wpclm = 1.479182934e-12 ppclm = -2.749357311e-19
+ pdiblc1 = 1.672174298e+00 lpdiblc1 = -2.367758932e-07 wpdiblc1 = -1.408078795e-11 ppdiblc1 = 2.617196056e-18
+ pdiblc2 = 4.684698606e-02 lpdiblc2 = -6.860232403e-09 wpdiblc2 = 2.059856486e-13 ppdiblc2 = -3.828655251e-20
+ pdiblcb = 9.254714851e-01 lpdiblcb = -1.968581093e-07 wpdiblcb = 4.377828398e-11 ppdiblcb = -8.137069644e-18
+ drout = -2.162511566e+00 ldrout = 4.929418876e-07 wdrout = 4.216895527e-11 pdrout = -7.837943716e-18
+ pscbe1 = 800000000.0
+ pscbe2 = -2.076171126e-09 lpscbe2 = 1.623203347e-15 wpscbe2 = -2.133815779e-19 ppscbe2 = 3.966123388e-26
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.459132804e+01 lbeta0 = -9.916237430e-07 wbeta0 = 2.568908610e-11 pbeta0 = -4.774830444e-18
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.395172510e-09 lagidl = 3.010800586e-16 wagidl = 3.595391044e-19 pagidl = -6.682753334e-26
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.934738292e-01 lkt1 = -2.693370996e-08 wkt1 = 1.016911632e-12 pkt1 = -1.890133641e-19
+ kt2 = 2.336833725e-01 lkt2 = -5.142806780e-08 wkt2 = 1.735882893e-12 pkt2 = -3.226485534e-19
+ at = 2.014816580e+05 lat = -2.793545395e-02 wat = -6.360928495e-07 pat = 1.182305780e-13
+ ute = -1.508684514e+00 lute = 2.343791916e-07 wute = -3.958932316e-12 pute = 7.358467498e-19
+ ua1 = -2.657626559e-09 lua1 = 5.301452092e-16 wua1 = -2.987467220e-20 pua1 = 5.552805322e-27
+ ub1 = 4.737798971e-18 lub1 = -8.121439041e-25 wub1 = 3.427805721e-29 pub1 = -6.371262494e-36
+ uc1 = -1.038108343e-10 luc1 = 1.276143166e-17 wuc1 = 2.399638041e-21 puc1 = -4.460207227e-28
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.81 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.098246063e+00 lvth0 = 7.294950629e-7
+ k1 = 4.276922968e-01 lk1 = 3.962872071e-7
+ k2 = 1.868581804e-02 lk2 = 5.621453833e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.092832443e-06 lcit = 2.417220556e-10 wcit = 1.694065895e-27 pcit = -5.421010862e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.791532993e-01 lvoff = 9.195555675e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.147437737e+00 lnfactor = -9.664292472e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.124081396e-02 lu0 = -3.340767752e-8
+ ua = -8.365019490e-10 lua = 3.589879299e-15
+ ub = 1.509438192e-18 lub = -9.691345396e-24
+ uc = -1.141297958e-10 luc = 8.465863493e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.012865143e+04 lvsat = 2.002511953e+0
+ a0 = 1.493812400e+00 la0 = -2.980908204e-6
+ ags = 1.038882350e-01 lags = 9.400718588e-7
+ a1 = 0.0
+ a2 = 1.012476349e+00 la2 = -4.247162113e-6
+ b0 = -1.285231938e-07 lb0 = 2.569033412e-12
+ b1 = 2.896927536e-09 lb1 = -5.790630792e-14
+ keta = 2.966561342e-02 lketa = -6.303652749e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.647222096e-02 lpclm = 3.146871810e-06 ppclm = -2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.516490733e-03 lpdiblc2 = -2.393052950e-8
+ pdiblcb = -2.424603954e-01 lpdiblcb = 1.745845204e-6
+ drout = 0.56
+ pscbe1 = 8.000121807e+08 lpscbe1 = -1.217936194e+0
+ pscbe2 = 1.121877068e-08 lpscbe2 = -1.158016781e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.498608750e-11 lalpha0 = 2.498330655e-15
+ alpha1 = -2.498608750e-11 lalpha1 = 2.498330655e-15
+ beta0 = 3.592705243e+01 lbeta0 = -5.926392753e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.263844868e-09 lagidl = -3.635470011e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.625313682e-02 legidl = 1.962312938e-5
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.376199758e-01 lkt1 = -6.299540746e-8
+ kt2 = -6.009202116e-02 lkt2 = 1.545849088e-7
+ at = 8.872762352e+04 lat = -1.773564932e+0
+ ute = -7.066532693e-02 lute = -1.231330245e-06 wute = 2.220446049e-22
+ ua1 = 2.157031712e-09 lua1 = -6.682427407e-15 wua1 = -6.617444900e-30
+ ub1 = -1.357081407e-18 lub1 = 1.281671407e-23
+ uc1 = -3.504300659e-11 luc1 = 5.253421821e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.82 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.061751
+ k1 = 0.44751769
+ k2 = 0.02149811
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.23314992
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1426029
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0095695
+ ua = -6.5690804e-10
+ ub = 1.02460111e-18
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.344684
+ ags = 0.150918
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.83 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-1
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595753e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 wpdiblc2 = -1.734723476e-24 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+3
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 wpscbe2 = -2.646977960e-29 ppscbe2 = -2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23 pub1 = -1.232595164e-44
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.84 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569066e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077653e-03 lketa = -3.715224604e-08 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = 4.440892099e-22 ppclm = -3.108624469e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048849e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807947e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123885e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.85 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-08 pk2 = -1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-06 pdsub = 1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = 5.898059818e-23 peta0 = 3.920475056e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = -9.367506770e-23 petab = -1.176142517e-27
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-9
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = 8.881784197e-22 pute = -2.220446049e-27
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.86 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.059631612e+00 lvth0 = 2.586054434e-8
+ k1 = 5.163379589e-01 lk1 = -1.485963682e-10
+ k2 = -3.690874683e-03 lk2 = -1.907482336e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.279561642e+00 ldsub = -4.971871951e-07 pdsub = 1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.986924020e-01 lvoff = -1.955441768e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.816966235e+00 lnfactor = 7.632892377e-7
+ eta0 = -4.398980000e-02 leta0 = 2.610515935e-07 peta0 = -4.440892099e-28
+ etab = -1.632772774e+00 letab = 7.979080824e-7
+ u0 = 8.012298384e-03 lu0 = 8.686250060e-10
+ ua = -7.759682813e-10 lua = 1.274097302e-16
+ ub = 6.727035311e-19 lub = 1.823100696e-25
+ uc = -9.895092236e-11 luc = 3.384048354e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.003651958e+04 lvsat = -2.626952517e-3
+ a0 = 1.678264962e+00 la0 = -4.701829257e-7
+ ags = -3.625107542e-01 lags = 7.883081324e-7
+ a1 = 0.0
+ a2 = 1.009669841e+00 la2 = -9.572104471e-9
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.793248020e-03 lketa = -2.322682382e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.567025060e+00 lpclm = -7.524585059e-7
+ pdiblc1 = 6.637643939e-02 lpdiblc1 = -2.707173962e-8
+ pdiblc2 = 8.111861681e-04 lpdiblc2 = -3.769435660e-10
+ pdiblcb = -3.034907083e-02 lpdiblcb = 5.289535676e-9
+ drout = 1.0
+ pscbe1 = 7.729094317e+08 lpscbe1 = 1.324376613e+1
+ pscbe2 = 9.028731239e-09 lpscbe2 = 1.463768495e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.609000049e+00 lbeta0 = 1.047440030e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.165212580e-10 lagidl = -3.050311102e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.213729371e-01 lkt1 = -5.704969315e-8
+ kt2 = -6.409955753e-02 lkt2 = 1.536741214e-8
+ at = 8.783879526e+04 lat = -2.578681467e-2
+ ute = -1.878857286e+00 lute = 8.214518228e-7
+ ua1 = -3.360596897e-09 lua1 = 2.897579860e-15 pua1 = -1.654361225e-36
+ ub1 = 4.154167712e-18 lub1 = -3.223006351e-24
+ uc1 = 3.233299061e-10 luc1 = -2.535572683e-16 wuc1 = -4.135903063e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.87 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.006613565e+00 lvth0 = -5.838818845e-11
+ k1 = 4.966170030e-01 lk1 = 9.492387336e-9
+ k2 = -1.761857806e-02 lk2 = 6.618088114e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.644100980e-01 ldsub = 2.576142694e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.427270611e-01 lvoff = 1.972806098e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.581462661e+00 lnfactor = -9.932013026e-8
+ eta0 = 0.49
+ etab = -1.216203250e-03 letab = 2.890215328e-10
+ u0 = 1.119413334e-02 lu0 = -6.868786489e-10
+ ua = -6.998804391e-11 lua = -2.177228284e-16
+ ub = 4.443627388e-19 lub = 2.939390328e-25
+ uc = -5.818012563e-11 luc = 1.390886414e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.048266764e+04 lvsat = 1.182103908e-2
+ a0 = 8.343866772e-01 la0 = -5.763614858e-8
+ ags = 9.847587520e-01 lags = 1.296684889e-7
+ a1 = 0.0
+ a2 = 1.171716763e+00 la2 = -8.879198318e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.192784488e-02 lketa = 2.058066866e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.557003024e-01 lpclm = 2.852782422e-07 wpclm = -4.440892099e-22 ppclm = -8.326672685e-29
+ pdiblc1 = -3.690848156e-01 lpdiblc1 = 1.858122041e-07 wpdiblc1 = -2.775557562e-22 ppdiblc1 = -2.775557562e-29
+ pdiblc2 = -8.705633412e-03 lpdiblc2 = 4.275544022e-09 wpdiblc2 = -6.722053469e-24 ppdiblc2 = 1.463672933e-30
+ pdiblcb = 1.686604462e-01 lpdiblcb = -9.200024691e-08 wpdiblcb = -1.110223025e-22
+ drout = 1.488187677e+00 ldrout = -2.386603096e-7
+ pscbe1 = 8.000276611e+08 lpscbe1 = -1.352270445e-2
+ pscbe2 = 9.493699522e-09 lpscbe2 = -8.093219498e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.555599215e+00 lbeta0 = 9.580609553e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.810185489e-10 lagidl = -4.323990079e-17
+ bgidl = 7.512236789e+08 lbgidl = 1.216192801e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.578143445e-01 lkt1 = 9.652417683e-9
+ kt2 = -1.325100891e-02 lkt2 = -9.490917822e-9
+ at = -2.296195638e+02 lat = 1.726719129e-2
+ ute = 4.373883268e-01 lute = -3.108911698e-07 pute = -2.220446049e-28
+ ua1 = 4.741250820e-09 lua1 = -1.063170433e-15
+ ub1 = -4.602396930e-18 lub1 = 1.057815405e-24
+ uc1 = -2.829276611e-10 luc1 = 4.282386859e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.88 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.786905057e-01 lvth0 = -5.450236936e-8
+ k1 = -4.472461707e-01 lk1 = 2.349529836e-7
+ k2 = 3.484937124e-01 lk2 = -8.083515471e-08 wk2 = 4.440892099e-22 pk2 = -5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.654947035e-01 ldsub = 1.071489094e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.427241235e-02 lvoff = -6.419405813e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.645192181e+00 lnfactor = -1.145432006e-7
+ eta0 = 6.885077223e-01 leta0 = -4.741753964e-8
+ etab = -6.25e-6
+ u0 = 1.813911423e-02 lu0 = -2.345826234e-9
+ ua = 1.276324974e-09 lua = -5.393166190e-16
+ ub = 9.196567555e-19 lub = 1.804055510e-25
+ uc = 2.387749767e-11 luc = -5.692240336e-18 wuc = 1.494418099e-32 puc = 4.543838814e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.449572143e+04 lvsat = 1.086244092e-2
+ a0 = -1.848840900e-01 la0 = 1.858370596e-7
+ ags = 2.197290171e+00 lags = -1.599688912e-7
+ a1 = 0.0
+ a2 = 1.355998444e+00 la2 = -1.328113483e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.115381286e-03 lketa = -1.013462857e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.298994868e-01 lpclm = 2.596102059e-8
+ pdiblc1 = 4.341255753e-01 lpdiblc1 = -6.050661960e-9
+ pdiblc2 = 7.396602975e-03 lpdiblc2 = 4.292028164e-10
+ pdiblcb = -4.163368351e-01 lpdiblcb = 4.773805368e-8
+ drout = 4.878551563e-01 ldrout = 2.891195681e-10
+ pscbe1 = 7.999012102e+08 lpscbe1 = 1.668263473e-2
+ pscbe2 = 1.518126485e-08 lpscbe2 = -1.439520925e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.233894147e+00 lbeta0 = 1.726517851e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.007565774e-10 lagidl = 7.184172364e-17
+ bgidl = 1.888486861e+09 lbgidl = -1.500387762e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.668066312e-01 lkt1 = -1.208659480e-8
+ kt2 = -7.705617102e-02 lkt2 = 5.750221250e-9
+ at = 1.224080320e+05 lat = -1.202726455e-2
+ ute = -2.351187446e+00 lute = 3.552159249e-7
+ ua1 = 5.215479907e-10 lua1 = -5.521001849e-17
+ ub1 = -1.482392574e-18 lub1 = 3.125399646e-25 wub1 = -1.540743956e-39
+ uc1 = -2.688967816e-10 luc1 = 3.947231239e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.89 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -2.062164096e-01 lvth0 = -1.663948370e-07 wvth0 = -7.740982042e-07 pvth0 = 1.438816332e-13
+ k1 = 1.181107242e+00 lk1 = -4.405654723e-08 wk1 = -9.754927563e-07 pk1 = 1.813148386e-13
+ k2 = -1.189255777e+00 lk2 = 1.968487362e-07 wk2 = 1.486384795e-06 pk2 = -2.762743418e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.828906208e+00 ldsub = -7.116787968e-07 wdsub = -2.145993095e-07 pdsub = 3.988757366e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 6.172330076e-02 lvoff = -7.575871627e-08 wvoff = -2.933987268e-07 pvoff = 5.453402136e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.905680794e+00 lnfactor = -9.179711862e-07 wnfactor = -7.499783272e-06 pnfactor = 1.393984717e-12
+ eta0 = 1.982978792e+00 leta0 = -2.927943610e-07 weta0 = -5.289517632e-07 peta0 = 9.831626422e-14
+ etab = -3.906706378e-01 letab = 7.261278975e-08 wetab = 4.713119458e-07 petab = -8.760275136e-14
+ u0 = 9.177474599e-04 lu0 = 6.189568656e-10 wu0 = 5.169917135e-09 pu0 = -9.609324978e-16
+ ua = 2.563693257e-09 lua = -8.328923095e-16 wua = -4.468017855e-15 pua = 8.304704788e-22
+ ub = 2.868112101e-18 lub = -1.635925700e-25 wub = -1.054397535e-25 pub = 1.959808699e-32
+ uc = -5.900652882e-11 luc = 9.140380651e-18 wuc = -2.074146127e-18 puc = 3.855215405e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.129705113e+06 lvsat = -1.934693159e-01 wvsat = -8.880794654e-01 pvsat = 1.650673302e-7
+ a0 = 7.135228311e+00 la0 = -1.156044173e-06 wa0 = -6.510018548e-06 pa0 = 1.210017148e-12
+ ags = 1.250000027e+00 lags = -5.081997045e-15 wags = -2.858905646e-14 pags = 5.313847140e-21
+ a1 = 0.0
+ a2 = -5.264002574e+00 la2 = 1.084278235e-06 wa2 = 4.812219417e-06 pa2 = -8.944472230e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.753488950e-01 lketa = 4.171850199e-08 wketa = -3.899072461e-08 pketa = 7.247205984e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.983923887e-01 lpclm = -5.850428111e-08 wpclm = 4.482155003e-09 ppclm = -8.330981505e-16
+ pdiblc1 = 2.089114339e+00 lpdiblc1 = -3.142725385e-07 wpdiblc1 = -4.359757601e-07 ppdiblc1 = 8.103481453e-14
+ pdiblc2 = 7.608195777e-02 lpdiblc2 = -1.229413660e-08 wpdiblc2 = -3.056852360e-08 ppdiblc2 = 5.681771482e-15
+ pdiblcb = -2.781768759e-01 lpdiblcb = 2.686401152e-08 wpdiblcb = 1.258604985e-06 ppdiblcb = -2.339369085e-13
+ drout = -2.162471648e+00 ldrout = 4.929344682e-07 wdrout = 4.305617551e-13 pdrout = -8.002851359e-20
+ pscbe1 = 7.999999958e+08 lpscbe1 = 7.849140167e-07 wpscbe1 = 4.415588379e-06 ppscbe1 = -8.207244873e-13
+ pscbe2 = -2.945237074e-08 lpscbe2 = 6.711617569e-15 wpscbe2 = 2.862494321e-14 ppscbe2 = -5.320518195e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.807219121e+01 lbeta0 = -1.638611781e-06 wbeta0 = -3.639641424e-06 pbeta0 = 6.765001515e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.724344829e-08 lagidl = 8.822899079e-15 wagidl = 4.794032536e-14 pagidl = -8.910668275e-21
+ bgidl = 9.999999970e+08 lbgidl = 5.590915680e-07 wbgidl = 3.145202637e-06 pbgidl = -5.845985413e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 4.692890577e-01 lkt1 = -1.872954478e-07 wkt1 = -9.021228384e-07 pkt1 = 1.676775720e-13
+ kt2 = 2.336850272e-01 lkt2 = -5.142837536e-08 wkt2 = 5.668548297e-15 pkt2 = -1.053613197e-21
+ at = 7.435873295e+05 lat = -1.286966351e-01 wat = -5.668382525e-01 pat = 1.053582260e-7
+ ute = -2.792624130e+00 lute = 4.730250480e-07 wute = 1.342511550e-06 pute = -2.495326218e-13
+ ua1 = -2.657655258e-09 lua1 = 5.301505435e-16 wua1 = 1.340311451e-22 pua1 = -2.491237098e-29
+ ub1 = 4.737832458e-18 lub1 = -8.121501283e-25 wub1 = -7.363307315e-31 pub1 = 1.368617919e-37
+ uc1 = -1.038085303e-10 luc1 = 1.276100342e-17 wuc1 = -9.410079440e-24 puc1 = 1.749051382e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.90 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.180836102e+00 lvth0 = 8.987579786e-06 wvth0 = 8.140255992e-08 pvth0 = -8.139349981e-12
+ k1 = 3.828265016e-01 lk1 = 4.882367371e-06 wk1 = 4.422071480e-08 pk1 = -4.421579303e-12
+ k2 = 1.232146936e-02 lk2 = 6.925785712e-07 wk2 = 6.272842076e-09 pk2 = -6.272143908e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.945947978e-05 lcit = 2.978082199e-09 wcit = 2.697316969e-11 pcit = -2.697016757e-15
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -3.832611055e-01 lvoff = 1.132917747e-05 wvoff = 1.026109442e-07 pvoff = -1.025995236e-11
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.158379199e+00 lnfactor = -1.190667409e-06 wnfactor = -1.078414628e-08 pnfactor = 1.078294601e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.502307589e-02 lu0 = -4.115917741e-07 wu0 = -3.727880570e-09 pu0 = 3.727465657e-13
+ ua = -1.242931393e-09 lua = 4.422830018e-14 wua = 4.005858019e-16 pua = -4.005412167e-20
+ ub = 2.606647261e-18 lub = -1.194000404e-22 wub = -1.081433397e-24 pub = 1.081313034e-28
+ uc = -2.099763664e-10 luc = 1.043017664e-14 wuc = 9.446848859e-17 puc = -9.445797425e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.665864420e+05 lvsat = 2.467149795e+01 wvsat = 2.234553838e-01 pvsat = -2.234305132e-5
+ a0 = 1.831296968e+00 la0 = -3.672560882e-05 wa0 = -3.326322151e-07 pa0 = 3.325951932e-11
+ ags = -2.542330341e-03 lags = 1.158194382e-05 wags = 1.049003067e-07 pags = -1.048886313e-11
+ a1 = 0.0
+ a2 = 1.493320298e+00 la2 = -5.232620520e-05 wa2 = -4.739303745e-07 pa2 = 4.738776261e-11
+ b0 = -4.193772130e-07 lb0 = 3.165119812e-11 wb0 = 2.866721201e-13 pb0 = -2.866402135e-17
+ b1 = 9.452810505e-09 lb1 = -7.134216378e-13 wb1 = -6.461622483e-15 pb1 = 6.460903305e-19
+ keta = 1.010326392e-01 lketa = -7.766273537e-06 wketa = -7.034091067e-08 pketa = 7.033308173e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.727464170e-01 lpclm = 3.877032609e-05 wpclm = 3.511516857e-07 ppclm = -3.511126025e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 4.225794026e-03 lpdiblc2 = -2.948307043e-07 wpdiblc2 = -2.670348931e-09 ppdiblc2 = 2.670051721e-13
+ pdiblcb = -4.401168727e-01 lpdiblcb = 2.150929302e-05 wpdiblcb = 1.948145725e-07 ppdiblcb = -1.947928896e-11
+ drout = 0.56
+ pscbe1 = 8.001500698e+08 lpscbe1 = -1.500530885e+01 wpscbe1 = -1.359065045e-01 ppscbe1 = 1.358913781e-5
+ pscbe2 = 2.432929831e-08 lpscbe2 = -1.426708520e-12 wpscbe2 = -1.292202446e-14 ppscbe2 = 1.292058623e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.078354692e-10 lalpha0 = 3.078012071e-14 walpha0 = 2.787825733e-16 palpha0 = -2.787515448e-20
+ alpha1 = -3.078354692e-10 lalpha1 = 3.078012071e-14 walpha1 = 2.787825733e-16 palpha1 = -2.787515448e-20
+ beta0 = 1.030229159e+02 lbeta0 = -7.301478847e-03 wbeta0 = -6.613115916e-05 pbeta0 = 6.612379877e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.379754997e-09 lagidl = -4.478999029e-13 wagidl = -4.056731573e-15 pagidl = 4.056280059e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -2.317892615e+00 legidl = 2.417623504e-04 wegidl = 2.189696746e-06 pegidl = -2.189453033e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.304879286e-01 lkt1 = -7.761207437e-07 wkt1 = -7.029502585e-09 pkt1 = 7.028720201e-13
+ kt2 = -7.759340585e-02 lkt2 = 1.904528587e-06 wkt2 = 1.724974978e-08 pkt2 = -1.724782988e-12
+ at = 2.895223996e+05 lat = -2.185080769e+01 wat = -1.979077488e-01 pat = 1.978857216e-5
+ ute = 6.874015874e-02 lute = -1.517032723e-05 wute = -1.374011136e-07 pute = 1.373858209e-11
+ ua1 = 2.913585076e-09 lua1 = -8.232934333e-14 wua1 = -7.456756393e-16 pua1 = 7.455926456e-20
+ ub1 = -2.808130188e-18 lub1 = 1.579054420e-22 wub1 = 1.430185601e-24 pub1 = -1.430026422e-28
+ uc1 = -9.451980607e-11 luc1 = 6.472360153e-15 wuc1 = 5.862164205e-17 puc1 = -5.861511747e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.91 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -5.111507366e-01 lvth0 = -4.398673926e-06 wvth0 = -5.426837328e-07 pvth0 = 4.335429792e-12
+ k1 = 7.466229913e-01 lk1 = -2.389513369e-06 wk1 = -2.948047653e-07 pk1 = 2.355156945e-12
+ k2 = 6.392710121e-02 lk2 = -3.389596950e-07 wk2 = -4.181894717e-08 pk2 = 3.340861325e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.924443156e-04 lcit = -1.457523920e-09 wcit = -1.798211312e-10 pcit = 1.436567641e-15
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 4.609021214e-01 lvoff = -5.544691532e-06 wvoff = -6.840729612e-07 pvoff = 5.464969957e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.069659816e+00 lnfactor = 5.827328171e-07 wnfactor = 7.189430854e-08 pnfactor = -5.743542847e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = -1.564557954e-02 lu0 = 2.014399925e-07 wu0 = 2.485253713e-08 pu0 = -1.985436883e-13
+ ua = 2.052621590e-09 lua = -2.164607997e-14 wua = -2.670572013e-15 pua = 2.133485263e-20
+ ub = -6.290126019e-18 lub = 5.843640412e-23 wub = 7.209555982e-24 pub = -5.759620550e-29
+ uc = 5.672002282e-10 luc = -5.104705282e-15 wuc = -6.297899239e-16 puc = 5.031309830e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.671743956e+06 lvsat = -1.207464939e+01 wvsat = -1.489702558e+00 pvsat = 1.190104008e-5
+ a0 = -9.052131216e-01 la0 = 1.797413562e-05 wa0 = 2.217548101e-06 pa0 = -1.771570350e-11
+ ags = 8.604551022e-01 lags = -5.668399670e-06 wags = -6.993353778e-07 pags = 5.586899420e-12
+ a1 = 0.0
+ a2 = -2.405626326e+00 la2 = 2.560933198e-05 wa2 = 3.159535830e-06 pa2 = -2.524112101e-11
+ b0 = 1.939026795e-06 lb0 = -1.549063299e-11 wb0 = -1.911147467e-12 pb0 = 1.526790867e-17
+ b1 = -4.370588646e-08 lb1 = 3.491606451e-13 wb1 = 4.307748322e-14 pb1 = -3.441404134e-19
+ keta = -4.776503718e-01 lketa = 3.800945941e-06 wketa = 4.689394045e-07 pketa = -3.746295940e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.516120287e+00 lpclm = -1.897485491e-05 wpclm = -2.341011238e-06 ppclm = 1.870203445e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.774272394e-02 lpdiblc2 = 1.442951454e-07 wpdiblc2 = 1.780232621e-08 ppdiblc2 = -1.422204698e-13
+ pdiblcb = 1.162590319e+00 lpdiblcb = -1.052701268e-05 wpdiblcb = -1.298763817e-06 ppdiblcb = 1.037565529e-11
+ drout = 0.56
+ pscbe1 = 7.990319895e+08 lpscbe1 = 7.343852554e+00 wpscbe1 = 9.060433631e-01 ppscbe1 = -7.238262642e-6
+ pscbe2 = -8.197805468e-08 lpscbe2 = 6.982553387e-13 wpscbe2 = 8.614682971e-14 ppscbe2 = -6.882158234e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.985662544e-09 lalpha0 = -1.506431293e-14 walpha0 = -1.858550488e-15 palpha0 = 1.484771824e-20
+ alpha1 = 1.985662544e-09 lalpha1 = -1.506431293e-14 walpha1 = -1.858550488e-15 palpha1 = 1.484771824e-20
+ beta0 = -4.410271673e+02 lbeta0 = 3.573467540e-03 wbeta0 = 4.408743944e-04 pbeta0 = -3.522088223e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.699430313e-08 lagidl = 2.192098063e-13 wagidl = 2.704487715e-14 pagidl = -2.160580078e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.569637951e+01 legidl = -1.183225932e-04 wegidl = -1.459797831e-05 pegidl = 1.166213510e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.883184811e-01 lkt1 = 3.798466506e-07 wkt1 = 4.686335057e-08 pkt1 = -3.743852154e-13
+ kt2 = 6.431742593e-02 lkt2 = -9.321085807e-07 wkt2 = -1.149983319e-07 pkt2 = 9.187067235e-13
+ at = -1.338631840e+06 lat = 1.069415575e+01 wat = 1.319384992e+00 pat = -1.054039518e-5
+ ute = -1.061636024e+00 lute = 7.424615349e-06 wute = 9.160074240e-07 pute = -7.317864229e-12
+ ua1 = -3.220964791e-09 lua1 = 4.029337646e-14 wua1 = 4.971170929e-15 pua1 = -3.971403830e-20
+ ub1 = 8.957769659e-18 lub1 = -7.728160049e-23 wub1 = -9.534570676e-24 pub1 = 7.617044564e-29
+ uc1 = 3.877507248e-10 luc1 = -3.167682794e-15 wuc1 = -3.908109470e-16 puc1 = 3.122137850e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.92 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16 wua = -1.654361225e-30
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-1
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595752e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 wpdiblc2 = 8.673617380e-25
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+3
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15 wagidl = -1.654361225e-30
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23 pub1 = 1.232595164e-44
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.93 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569065e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077653e-03 lketa = -3.715224604e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = 3.330669074e-22 ppclm = 2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048848e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807946e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123885e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.94 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = 5.377642776e-23 peta0 = -2.185751580e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = 3.920475056e-22 petab = 4.631711681e-28
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-9
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16 pagidl = 4.135903063e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-02 wat = 2.328306437e-16
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = -4.440892099e-22 pute = -6.661338148e-28
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24 pub1 = 6.162975822e-45
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.95 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.047616465e+00 lvth0 = 1.397912612e-08 wvth0 = -1.184239303e-08 pvth0 = 1.171058719e-14
+ k1 = 4.467500259e-01 lk1 = 6.866482286e-08 wk1 = 6.858739762e-08 pk1 = -6.782401988e-14
+ k2 = 3.540557254e-02 lk2 = -3.885205200e-08 wk2 = -3.853431850e-08 pk2 = 3.810543154e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.912433260e+00 ldsub = -1.123014953e-06 wdsub = -6.237721905e-07 pdsub = 6.168296060e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.426527285e-01 lvoff = -3.571003769e-07 wvoff = -3.364372703e-07 pvoff = 3.326927234e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.256158503e+01 lnfactor = 1.498180722e-05 wnfactor = 1.417181645e-05 pnfactor = -1.401408413e-11
+ eta0 = -4.574898055e-01 leta0 = 6.699493440e-07 weta0 = 4.075547024e-07 peta0 = -4.030186186e-13
+ etab = -1.633094605e+00 letab = 7.982263309e-07 wetab = 3.172031693e-10 petab = -3.136726980e-16
+ u0 = -3.130665353e-02 lu0 = 3.974995698e-08 wu0 = 3.875362402e-08 pu0 = -3.832229619e-14
+ ua = -8.360635370e-09 lua = 7.627659475e-15 wua = 7.475614746e-15 pua = -7.392411154e-21
+ ub = 2.781703904e-18 lub = -1.903217129e-24 wub = -2.078677165e-24 pub = 2.055541488e-30
+ uc = -1.149161555e-10 luc = 4.962802368e-17 wuc = 1.573568506e-17 puc = -1.556054688e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.749760186e+05 lvsat = -4.228368749e-01 wvsat = -4.188297189e-01 pvsat = 4.141681441e-7
+ a0 = 2.019660525e+00 la0 = -8.077787556e-07 wa0 = -3.364869772e-07 pa0 = 3.327418771e-13
+ ags = -3.625107549e-01 lags = 7.883081331e-07 wags = 6.444036416e-16 pags = -6.372316008e-22
+ a1 = 0.0
+ a2 = 5.823493325e-01 la2 = 4.129923269e-07 wa2 = 4.211764944e-07 pa2 = -4.164888000e-13
+ b0 = 9.707705920e-16 lb0 = -9.599659153e-22 wb0 = -9.568128524e-22 pb0 = 9.461635254e-28
+ b1 = 4.035937759e-19 lb1 = -3.991017772e-25 wb1 = -3.977909046e-25 pb1 = 3.933634918e-31
+ keta = 4.804604229e-03 lketa = -1.829370363e-08 wketa = 4.916917070e-09 pketa = -4.862191783e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.914299633e+00 lpclm = -1.095867913e-06 wpclm = -3.422814592e-07 ppclm = 3.384718665e-13
+ pdiblc1 = 1.168996606e-01 lpdiblc1 = -7.703263734e-08 wpdiblc1 = -4.979679830e-08 ppdiblc1 = 4.924255993e-14
+ pdiblc2 = 1.466407932e-03 lpdiblc2 = -1.024872712e-09 wpdiblc2 = -6.458009852e-10 ppdiblc2 = 6.386132203e-16
+ pdiblcb = -2.066815844e-01 lpdiblcb = 1.796594684e-07 wpdiblcb = 1.737972047e-07 ppdiblcb = -1.718628418e-13
+ drout = 5.811830963e-01 ldrout = 4.141554715e-07 wdrout = 4.127951542e-07 pdrout = -4.082007441e-13
+ pscbe1 = 2.050336954e+08 lpscbe1 = 5.747990455e+02 wpscbe1 = 5.597108190e+02 ppscbe1 = -5.534812376e-4
+ pscbe2 = 6.811211336e-08 lpscbe2 = -5.827940723e-14 wpscbe2 = -5.823388125e-14 ppscbe2 = 5.758573815e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.343431244e+00 lbeta0 = 1.310053054e-06 wbeta0 = 2.617504563e-07 pbeta0 = -2.588371737e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.314897187e-09 lagidl = 1.802664647e-15 wagidl = 2.100772911e-15 pagidl = -2.077391308e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.748677571e-01 lkt1 = -1.030372705e-07 wkt1 = -4.583652852e-08 pkt1 = 4.532636795e-14
+ kt2 = -8.716677806e-02 lkt2 = 3.817789451e-08 wkt2 = 2.273556004e-08 pkt2 = -2.248251325e-14
+ at = 1.263791376e+05 lat = -6.389820300e-02 wat = -3.798620930e-02 pat = 3.756342279e-8
+ ute = -1.913227686e+00 lute = 8.554396804e-07 wute = 3.387622248e-08 pute = -3.349918012e-14
+ ua1 = -4.133738016e-09 lua1 = 3.662115918e-15 wua1 = 7.620248955e-16 pua1 = -7.535435584e-22
+ ub1 = 5.503375746e-18 lub1 = -4.557197700e-24 wub1 = -1.329809122e-24 pub1 = 1.315008346e-30
+ uc1 = 4.331615978e-10 luc1 = -3.621665333e-16 wuc1 = -1.082525317e-16 puc1 = 1.070476810e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.96 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.297338687e+00 lvth0 = 1.360608290e-07 wvth0 = 2.865450765e-07 pvth0 = -1.341620951e-13
+ k1 = 1.084757674e+00 lk1 = -2.432379762e-07 wk1 = -5.796843847e-07 pk1 = 2.490966063e-13
+ k2 = -3.452969821e-01 lk2 = 1.472620059e-07 wk2 = 3.229670439e-07 pk2 = -1.386217395e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.848905686e+00 ldsub = 7.157908182e-07 wdsub = 1.561713711e-06 pdsub = -4.515888864e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.065666696e+00 lvoff = 2.336107399e-07 wvoff = 8.111074084e-07 pvoff = -2.283074436e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.300137660e+01 lnfactor = -7.292557829e-06 wnfactor = -2.899691442e-05 pnfactor = 7.089813327e-12
+ eta0 = 1.317000017e+00 leta0 = -1.975454955e-07 weta0 = -8.151094106e-07 peta0 = 1.947051863e-13
+ etab = -1.281599537e-03 letab = 4.819070393e-10 wetab = 6.445601891e-11 petab = -1.901121986e-16
+ u0 = 8.594045236e-02 lu0 = -1.756863567e-08 wu0 = -7.367161644e-08 pu0 = 1.663903112e-14
+ ua = 1.420332019e-08 lua = -3.403181479e-15 wua = -1.406808661e-14 pua = 3.139658126e-21
+ ub = -3.440248070e-18 lub = 1.138508533e-24 wub = 3.828757875e-24 pub = -8.324262797e-31
+ uc = -3.747081394e-11 luc = 1.176731953e-17 wuc = -2.041155320e-17 puc = 2.110753484e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.476545150e+05 lvsat = 1.748705140e-01 wvsat = 7.570929062e-01 pvsat = -1.607051496e-7
+ a0 = 3.949277881e-01 la0 = -1.349566276e-08 wa0 = 4.331403492e-07 pa0 = -4.350583392e-14
+ ags = 7.469353827e-01 lags = 2.459331998e-07 wags = 2.344039449e-07 pags = -1.145930569e-13
+ a1 = 0.0
+ a2 = 1.983329918e+00 la2 = -2.719050519e-07 wa2 = -7.999437809e-07 pa2 = 1.804802690e-13
+ b0 = -1.941541184e-15 lb0 = 4.637759426e-22 wb0 = 1.913625705e-21 pb0 = -4.571077721e-28
+ b1 = -8.071875518e-19 lb1 = 1.928128905e-25 wb1 = 7.955818092e-25 pb1 = -1.900406268e-31
+ keta = -1.416863263e-02 lketa = -9.018257333e-09 wketa = -2.736009030e-08 pketa = 1.091706881e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.265185887e+00 lpclm = 4.584871736e-07 wpclm = 6.992846010e-07 ppclm = -1.707185333e-13
+ pdiblc1 = -5.151856770e-01 lpdiblc1 = 2.319749217e-07 wpdiblc1 = 1.440002233e-07 ppdiblc1 = -4.549899001e-14
+ pdiblc2 = -1.668860894e-02 lpdiblc2 = 7.850570385e-09 wpdiblc2 = 7.868196303e-09 ppdiblc2 = -3.523624634e-15
+ pdiblcb = -2.523915908e-01 lpdiblcb = 2.020057192e-07 wpdiblcb = 4.149981508e-07 ppdiblcb = -2.897787484e-13
+ drout = 2.754316326e+00 ldrout = -6.482241706e-07 wdrout = -1.247924252e-06 pdrout = 4.036751518e-13
+ pscbe1 = 1.935803422e+09 lpscbe1 = -2.713223510e+02 wpscbe1 = -1.119445577e+03 ppscbe1 = 2.674079500e-4
+ pscbe2 = -1.120279352e-07 lpscbe2 = 2.978565831e-14 wpscbe2 = 1.197743967e-13 ppscbe2 = -2.943716867e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.581254503e+00 lbeta0 = 2.160483970e-07 wbeta0 = -2.528641655e-08 pbeta0 = -1.185134577e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.479120858e-09 lagidl = -5.409869541e-16 wagidl = -3.152119994e-15 pagidl = 4.905904462e-22
+ bgidl = 5.281633166e+08 lbgidl = 2.306667994e+02 wbgidl = 2.198532004e+02 pbgidl = -1.074796341e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.101814353e-01 lkt1 = 6.088752738e-08 wkt1 = 1.501763568e-07 pkt1 = -5.049845129e-14
+ kt2 = 3.472639696e-02 lkt2 = -2.141202197e-08 wkt2 = -4.728758674e-08 pkt2 = 1.174970251e-14
+ at = -1.224106452e+05 lat = 5.772765811e-02 wat = 1.204243068e-01 pat = -3.987872624e-8
+ ute = 8.255450053e-01 lute = -4.834641252e-07 wute = -3.825757618e-07 pute = 1.700917015e-13
+ ua1 = 6.337484800e-09 lua1 = -1.456950780e-15 wua1 = -1.573283328e-15 pua1 = 3.881185728e-22
+ ub1 = -7.250399985e-18 lub1 = 1.677740641e-24 wub1 = 2.609930067e-24 pub1 = -6.110119511e-31
+ uc1 = -4.402376540e-10 luc1 = 6.481215895e-17 wuc1 = 1.550481898e-16 puc1 = -2.167214271e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.97 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -6.176616124e-01 lvth0 = -2.629363391e-08 wvth0 = -1.587136199e-07 pvth0 = -2.780315025e-14
+ k1 = 2.500047514e+00 lk1 = -5.813082601e-07 wk1 = -2.904917496e-06 pk1 = 8.045250396e-13
+ k2 = -1.157335456e+00 lk2 = 3.412336362e-07 wk2 = 1.484178357e-06 pk2 = -4.160002858e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.734633138e+01 ldsub = 4.417660893e-06 wdsub = 1.745716545e-05 pdsub = -4.248535442e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.341235372e-01 lvoff = -5.298315299e-08 wvoff = -9.841546538e-08 pvoff = -1.104971475e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.983020398e+01 lnfactor = -4.146359823e-06 wnfactor = -1.595230370e-05 pnfactor = 3.973847163e-12
+ eta0 = -4.452025897e+00 leta0 = 1.180501725e-06 weta0 = 5.066623027e-06 peta0 = -1.210264241e-12
+ etab = -7.447189740e-01 letab = 1.780667927e-07 wetab = 7.340052444e-07 petab = -1.755065483e-13
+ u0 = 3.684682341e-02 lu0 = -5.841640523e-09 wu0 = -1.843872973e-08 pu0 = 3.445551471e-15
+ ua = 7.440939352e-09 lua = -1.787851569e-15 wua = -6.075979553e-15 pua = 1.230583514e-21
+ ub = -4.271439599e-18 lub = 1.337055253e-24 wub = 5.116458771e-24 pub = -1.140019393e-30
+ uc = 3.347570743e-10 luc = -7.714675613e-17 wuc = -3.064097501e-16 puc = 7.042714277e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.133665286e+06 lvsat = 2.670769070e-01 wvsat = 1.141508969e+00 pvsat = -2.525306145e-7
+ a0 = 4.891591352e+00 la0 = -1.087613688e-06 wa0 = -5.003485878e-06 pa0 = 1.255141073e-12
+ ags = 3.046659586e+00 lags = -3.034019207e-07 wags = -8.371571814e-07 pags = 1.413707494e-13
+ a1 = 0.0
+ a2 = 3.576415423e+00 la2 = -6.524453865e-07 wa2 = -2.188491824e-06 pa2 = 5.121627400e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.356768448e+00 lketa = -3.364939978e-07 wketa = -1.328276511e-06 pketa = 3.216669743e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.097820927e+00 lpclm = 4.185087055e-07 wpclm = 1.604317049e-06 ppclm = -3.869036343e-13
+ pdiblc1 = -5.701544345e+00 lpdiblc1 = 1.470840417e-06 wpdiblc1 = 6.047451258e-06 ppdiblc1 = -1.455656339e-12
+ pdiblc2 = -1.347910092e-01 lpdiblc2 = 3.606169074e-08 wpdiblc2 = 1.401432387e-07 ppdiblc2 = -3.512016401e-14
+ pdiblcb = -4.372307801e+00 lpdiblcb = 1.186130104e-06 wpdiblcb = 3.899092016e-06 ppdiblcb = -1.122024250e-12
+ drout = 1.289711006e+01 ldrout = -3.071033310e-06 wdrout = -1.223083464e-05 pdrout = 3.027162956e-12
+ pscbe1 = 7.998144663e+08 lpscbe1 = 3.133096612e-02 wpscbe1 = 8.549668424e-02 ppscbe1 = -1.443771768e-8
+ pscbe2 = 4.686327011e-08 lpscbe2 = -8.168683898e-15 wpscbe2 = -3.122648139e-14 ppscbe2 = 6.632411069e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.467118439e+01 lbeta0 = 5.770358476e-06 wbeta0 = 2.257574932e-05 pbeta0 = -5.517222864e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.728238588e-09 lagidl = -6.004937064e-16 wagidl = -3.872504073e-15 pagidl = 6.626685912e-22
+ bgidl = 2.685132204e+09 lbgidl = -2.845683587e+02 wbgidl = -7.851911759e+02 pbgidl = 1.325953161e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.971956461e-01 lkt1 = -6.164938809e-08 wkt1 = -2.657345183e-07 pkt1 = 4.885017945e-14
+ kt2 = -1.537970646e+00 lkt2 = 3.542581206e-07 wkt2 = 1.439909446e-06 pkt2 = -3.434970528e-13
+ at = 1.238074386e+04 lat = 2.553003901e-02 wat = 1.084453158e-01 pat = -3.701730465e-8
+ ute = 1.907099889e+00 lute = -7.418151404e-07 wute = -4.197061680e-06 pute = 1.081257953e-12
+ ua1 = 1.533516198e-08 lua1 = -3.606225928e-15 wua1 = -1.460062385e-14 pua1 = 3.499959402e-21
+ ub1 = -2.462906326e-17 lub1 = 5.828981938e-24 wub1 = 2.281386785e-23 pub1 = -5.437126570e-30
+ uc1 = -1.307216976e-10 luc1 = -9.121917570e-18 wuc1 = -1.361884026e-16 puc1 = 4.789554212e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.98 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 7.331292215e-01 lvth0 = -2.800120841e-07 wvth0 = -1.699937924e-06 pvth0 = 2.558652915e-13
+ k1 = -1.049609291e+01 lk1 = 1.775764550e-06 wk1 = 1.053381261e-05 pk1 = -1.612340871e-12
+ k2 = 6.133871344e+00 lk2 = -9.796312703e-07 wk2 = -5.731450404e-06 pk2 = 8.832902352e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.324281792e+01 ldsub = -8.258022104e-06 wdsub = -4.793241580e-05 pdsub = 7.477729557e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.091684080e+00 lvoff = -2.362987002e-07 wvoff = -1.308550730e-06 pvoff = 2.127657614e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -3.974058775e+01 lnfactor = 6.508652701e-06 wnfactor = 3.946142723e-05 pnfactor = -5.925859172e-12
+ eta0 = 1.518504107e+01 leta0 = -2.350599804e-06 weta0 = -1.354119479e-05 peta0 = 2.126534580e-12
+ etab = 1.523527716e+00 letab = -2.256063863e-07 wetab = -1.415364064e-06 petab = 2.063286293e-13
+ u0 = 1.150529575e-02 lu0 = -1.719483787e-09 wu0 = -5.265403390e-09 pu0 = 1.343886055e-15
+ ua = -5.049960985e-09 lua = 3.538505724e-16 wua = 3.036167266e-15 pua = -3.392094139e-22
+ ub = 1.314208153e-17 lub = -1.764995698e-24 wub = -1.023169005e-23 pub = 1.597976241e-30
+ uc = -7.544714579e-10 luc = 1.175418525e-16 wuc = 6.833913882e-16 puc = -1.064573539e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.475830425e+06 lvsat = -3.769336546e-01 wvsat = -2.214850187e+00 pvsat = 3.458938186e-7
+ a0 = -8.134220272e+00 la0 = 1.224004769e-06 wa0 = 8.539885903e-06 pa0 = -1.135811450e-12
+ ags = 1.249999397e+00 lags = 9.398935319e-14 wags = 5.923722171e-13 pags = -9.233305676e-20
+ a1 = 0.0
+ a2 = -1.062188100e+01 la2 = 1.920910844e-06 wa2 = 1.009306226e-05 pa2 = -1.719050729e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.899529475e+00 lketa = 6.066195312e-07 wketa = 3.533081387e-06 pketa = -5.495316762e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.315703600e+00 lpclm = -7.314421811e-07 wpclm = -4.250754756e-06 ppclm = 6.624293007e-13
+ pdiblc1 = 1.826469387e+01 lpdiblc1 = -2.835696021e-06 wpdiblc1 = -1.637898281e-05 ppdiblc1 = 2.566205270e-12
+ pdiblc2 = 5.027718896e-01 lpdiblc2 = -7.881182538e-08 wpdiblc2 = -4.511235076e-07 ppdiblc2 = 7.124306893e-14
+ pdiblcb = 1.696530174e+01 lpdiblcb = -2.660484668e-06 wpdiblcb = -1.573694690e-05 ppdiblcb = 2.414773072e-12
+ drout = -3.796252626e+01 ldrout = 6.073088969e-06 wdrout = 3.528532186e-05 pdrout = -5.499923119e-12
+ pscbe1 = 7.999999963e+08 lpscbe1 = 5.753192902e-07 wpscbe1 = 3.940093994e-06 ppscbe1 = -6.141414642e-13
+ pscbe2 = -8.034473494e-08 lpscbe2 = 1.465313350e-14 wpscbe2 = 7.878557700e-14 ppscbe2 = -1.314785101e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.157188191e+01 lbeta0 = -1.153744315e-05 wbeta0 = -6.622633357e-05 pbeta0 = 1.043300613e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.092969001e-09 lagidl = -1.711273415e-16 wagidl = 2.988890734e-16 pagidl = -4.595796661e-23
+ bgidl = 9.999969400e+08 lbgidl = 4.769605656e-04 wbgidl = 3.016208206e-03 pbgidl = -4.701363716e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 3.186927727e-01 lkt1 = -1.637437602e-07 wkt1 = -7.536918268e-07 pkt1 = 1.444645106e-13
+ kt2 = 3.968742406e+00 lkt2 = -6.336117692e-07 wkt2 = -3.681354719e-06 pkt2 = 5.738127599e-13
+ at = 1.445723757e+06 lat = -2.383153394e-01 wat = -1.258879362e+00 pat = 2.134008325e-7
+ ute = -1.667258710e+01 lute = 2.636913378e-06 wute = 1.502290841e-05 pute = -2.382308566e-12
+ ua1 = -4.116056328e-08 lua1 = 6.531598814e-15 wua1 = 3.794931334e-14 pua1 = -5.915159472e-21
+ ub1 = 6.372135967e-17 lub1 = -1.000591249e-23 wub1 = -5.813546279e-23 pub1 = 9.061574586e-30
+ uc1 = -1.030594110e-09 luc1 = 1.572190720e-16 wuc1 = 9.134602471e-16 puc1 = -1.423810487e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.99 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.100 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.110389418e+00 lvth0 = 3.885659956e-7
+ k1 = 4.210956021e-01 lk1 = 2.110826255e-7
+ k2 = 1.775005695e-02 lk2 = 2.994270855e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 pcit = 8.131516294e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.944604484e-01 lvoff = 4.898018407e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.149046479e+00 lnfactor = -5.147691352e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.179692641e-02 lu0 = -1.779462005e-8
+ ua = -8.962599665e-10 lua = 1.912151425e-15
+ ub = 1.670762721e-18 lub = -5.162101108e-24
+ uc = -1.282222813e-10 luc = 4.509347416e-16 wuc = 8.271806126e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.679434283e+04 lvsat = 1.066639228e+0
+ a0 = 1.543433334e+00 la0 = -1.587782595e-6
+ ags = 8.823956664e-02 lags = 5.007298559e-7
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = -1.712879585e-07 lb0 = 1.368397233e-12
+ b1 = 3.860850241e-09 lb1 = -3.084383066e-14
+ keta = 4.015882949e-02 lketa = -3.357644528e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 ppclm = -5.329070518e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.914844237e-03 lpdiblc2 = -1.274661131e-8
+ pdiblcb = -2.715221659e-01 lpdiblcb = 9.299255256e-07 wpdiblcb = 1.776356839e-21
+ drout = 0.56
+ pscbe1 = 8.000324548e+08 lpscbe1 = -6.487344657e-1
+ pscbe2 = 1.314643402e-08 lpscbe2 = -6.168183535e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.579227219e+01 lbeta0 = -3.156696758e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.869014186e-09 lagidl = -1.936435346e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.229045954e-01 legidl = 1.045227198e-05 wegidl = -1.776356839e-21
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365713387e-01 lkt1 = -3.355454267e-8
+ kt2 = -6.266527973e-02 lkt2 = 8.233974711e-8
+ at = 1.182508234e+05 lat = -9.446904559e-1
+ ute = -5.016829954e-02 lute = -6.558688149e-7
+ ua1 = 2.268269050e-09 lua1 = -3.559399084e-15
+ ub1 = -1.570431596e-18 lub1 = 6.826830664e-24
+ uc1 = -4.378798232e-11 luc1 = 2.798238376e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.101 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-01 pvsat = -7.450580597e-21
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595753e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 ppdiblc2 = -4.163336342e-29
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-07 wpdiblcb = 1.776356839e-21
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+03 wpscbe1 = 7.629394531e-12
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23 pub1 = -4.930380658e-44
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.102 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569065e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077654e-03 lketa = -3.715224604e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = -1.332267630e-21 ppclm = -4.440892099e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048848e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807946e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292611e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123884e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.103 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = -2.498001805e-22 peta0 = 9.922618283e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = -7.147060721e-22 petab = 7.910339050e-28
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-09 wu0 = 1.110223025e-22
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 pute = 1.776356839e-27
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24 pub1 = 2.465190329e-44
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.104 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.060692995e+00 lvth0 = 2.691011409e-8
+ k1 = 5.224851534e-01 lk1 = -6.227372655e-9
+ k2 = -7.144540537e-03 lk2 = 3.224478319e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.223655613e+00 ldsub = -4.419034005e-07 pdsub = -3.552713679e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.288458330e-01 lvoff = 1.026340558e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.087125419e+00 lnfactor = -4.927330750e-7
+ eta0 = -7.462418332e-03 leta0 = 2.249307616e-7
+ etab = -1.632744345e+00 letab = 7.978799692e-7
+ u0 = 1.148561965e-02 lu0 = -2.566038196e-9
+ ua = -1.059609635e-10 lua = -5.351404061e-16
+ ub = 4.864006036e-19 lub = 3.665394455e-25
+ uc = -9.754060033e-11 luc = 3.244585840e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.249860650e+04 lvsat = 3.449316359e-2
+ a0 = 1.648107076e+00 la0 = -4.403606970e-7
+ ags = -3.625107541e-01 lags = 7.883081323e-7
+ a1 = 0.0
+ a2 = 1.047418086e+00 la2 = -4.690021102e-8
+ b0 = -8.575503616e-17 lb0 = 8.480058261e-23
+ b1 = -3.565229431e-20 lb1 = 3.525548427e-26
+ keta = 1.023393023e-02 lketa = -2.366260124e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.536347840e+00 lpclm = -7.221227228e-7
+ pdiblc1 = 6.191336573e-02 lpdiblc1 = -2.265833997e-8
+ pdiblc2 = 7.533057929e-04 lpdiblc2 = -3.197073994e-10
+ pdiblcb = -1.477237207e-02 lpdiblcb = -1.011379443e-8
+ drout = 1.036997061e+00 ldrout = -3.658528362e-8
+ pscbe1 = 8.230739141e+08 lpscbe1 = -3.636238561e+1
+ pscbe2 = 3.809477986e-09 lpscbe2 = 5.307539814e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.632459620e+00 lbeta0 = 1.024241563e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.004804533e-09 lagidl = -4.912187918e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.254810687e-01 lkt1 = -5.298728500e-8
+ kt2 = -6.206186670e-02 lkt2 = 1.335240081e-08 wkt2 = -4.440892099e-22
+ at = 8.443425409e+04 lat = -2.242016604e-2
+ ute = -1.875821105e+00 lute = 8.184494349e-07 pute = -7.105427358e-27
+ ua1 = -3.292299871e-09 lua1 = 2.830042980e-15 wua1 = -6.617444900e-30 pua1 = 6.617444900e-36
+ ub1 = 4.034982618e-18 lub1 = -3.105147788e-24 pub1 = 1.232595164e-44
+ uc1 = 3.136276955e-10 luc1 = -2.439630433e-16 wuc1 = 8.271806126e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.105 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.809317576e-01 lvth0 = -1.208276190e-8
+ k1 = 4.446623754e-01 lk1 = 3.181784882e-8
+ k2 = 1.132757422e-02 lk2 = -5.805984424e-09 wk2 = -6.938893904e-24 pk2 = -1.040834086e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.244403898e-01 ldsub = 2.171402925e-07 pdsub = 8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.700309796e-01 lvoff = -1.848941181e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.825934693e-01 lnfactor = 5.361094594e-7
+ eta0 = 4.169452362e-01 leta0 = 1.745059157e-8
+ etab = -1.210426333e-03 letab = 2.719825911e-10
+ u0 = 4.591262030e-03 lu0 = 8.044064145e-10
+ ua = -1.330850367e-09 lua = 6.367127645e-17
+ ub = 7.875179014e-19 lub = 2.193322321e-25
+ uc = -6.000952568e-11 luc = 1.409804193e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.833766079e+04 lvsat = -2.582274881e-3
+ a0 = 8.732071908e-01 la0 = -6.153539006e-8
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 1.100021230e+00 la2 = -7.261631000e-8
+ b0 = 1.715100723e-16 lb0 = -4.096861098e-23
+ b1 = 7.130458861e-20 lb1 = -1.703252708e-26
+ keta = -4.438001254e-02 lketa = 3.036516966e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.930264200e-01 lpclm = 2.699774716e-07 wpclm = 1.776356839e-21
+ pdiblc1 = -3.561786926e-01 lpdiblc1 = 1.817343246e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = -5.551115123e-29
+ pdiblc2 = -8.000440691e-03 lpdiblc2 = 3.959736644e-09 wpdiblc2 = 6.071532166e-24 ppdiblc2 = -1.170938346e-29
+ pdiblcb = 2.058549522e-01 lpdiblcb = -1.179718745e-07 wpdiblcb = -4.440892099e-22 ppdiblcb = 4.440892099e-28
+ drout = 1.376341573e+00 ldrout = -2.024806355e-7
+ pscbe1 = 6.996965507e+08 lpscbe1 = 2.395310605e+1
+ pscbe2 = 2.022856548e-08 lpscbe2 = -2.719259489e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.553332902e+00 lbeta0 = 8.518424213e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.492459760e-12 lagidl = 7.296188029e-19
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.443546811e-01 lkt1 = 5.126457872e-9
+ kt2 = -1.748919269e-02 lkt2 = -8.437842332e-9
+ at = 1.056349506e+04 lat = 1.369303193e-2
+ ute = 4.030997005e-01 lute = -2.956465794e-07 wute = -1.776356839e-21
+ ua1 = 4.600244176e-09 lua1 = -1.028385029e-15
+ ub1 = -4.368480081e-18 lub1 = 1.003053022e-24
+ uc1 = -2.690313562e-10 luc1 = 4.088148730e-17 wuc1 = -1.654361225e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.106 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.929153274e-01 lvth0 = -5.699424658e-8
+ k1 = -7.076014787e-01 lk1 = 3.070591157e-7
+ k2 = 4.815142591e-01 lk2 = -1.181194778e-07 wk2 = -4.440892099e-22 pk2 = 2.775557562e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.930105641e+00 ldsub = -2.736291180e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 2.545185588e-02 lvoff = -6.518439671e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.215455554e+00 lnfactor = 2.416156933e-7
+ eta0 = 1.142607435e+00 leta0 = -1.558883378e-7
+ etab = 6.577949496e-02 letab = -1.572989991e-08 wetab = 2.220446049e-22 petab = 1.864827737e-29
+ u0 = 1.648652989e-02 lu0 = -2.037016219e-9
+ ua = 7.317609614e-10 lua = -4.290246915e-16
+ ub = 1.378223032e-18 lub = 7.823049762e-26
+ uc = -3.584695304e-12 luc = 6.198427007e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.268042791e+05 lvsat = -1.177079600e-2
+ a0 = -6.333250901e-01 la0 = 2.983299759e-7
+ ags = 2.122259360e+00 lags = -1.472984367e-7
+ a1 = 0.0
+ a2 = 1.159853299e+00 la2 = -8.690839645e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.099323509e-01 lketa = 1.869500404e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.736875497e-01 lpclm = -8.715494325e-9
+ pdiblc1 = 9.761327191e-01 lpdiblc1 = -1.365149023e-7
+ pdiblc2 = 1.995704097e-02 lpdiblc2 = -2.718466999e-9
+ pdiblcb = -6.687792477e-02 lpdiblcb = -5.282417213e-8
+ drout = -6.083421450e-01 ldrout = 2.716007644e-7
+ pscbe1 = 7.999088729e+08 lpscbe1 = 1.538864396e-2
+ pscbe2 = 1.238256912e-08 lpscbe2 = -8.450863393e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025726182e+01 lbeta0 = -3.218332598e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -5.478325244e-10 lagidl = 1.312338700e-16 wagidl = 2.326445473e-31 pagidl = 8.401053096e-38
+ bgidl = 1.818113540e+09 lbgidl = -1.381548262e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.906232774e-01 lkt1 = -7.708362526e-9
+ kt2 = 5.199674285e-02 lkt2 = -2.503594776e-8
+ at = 1.321275210e+05 lat = -1.534496695e-2
+ ute = -2.727352100e+00 lute = 4.521244422e-7
+ ua1 = -7.870433631e-10 lua1 = 2.584763459e-16 pua1 = -8.271806126e-37
+ ub1 = 5.623166473e-19 lub1 = -1.747663926e-25
+ uc1 = -2.811027645e-10 luc1 = 4.376498461e-17 wuc1 = 1.654361225e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.107 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.743799556e+00 lvth0 = 1.140090424e-07 wvth0 = 5.432232694e-07 pvth0 = -1.009689091e-13
+ k1 = 2.232319638e+00 lk1 = -2.084726409e-07 wk1 = -9.933178159e-07 pk1 = 1.846279824e-13
+ k2 = 8.272327637e-01 lk2 = -1.942691642e-07 wk2 = -9.256417598e-07 pk2 = 1.720490339e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.564914671e-01 ldsub = -4.586146319e-08 wdsub = -2.185194647e-07 pdsub = 4.061621291e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.926102424e-02 lvoff = -6.157697174e-08 wvoff = -2.933981828e-07 pvoff = 5.453392024e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.211461117e+01 lnfactor = -1.574017114e-06 wnfactor = -7.499781732e-06 pnfactor = 1.393984431e-12
+ eta0 = 8.167465371e-01 leta0 = -1.110137198e-07 weta0 = -5.289511586e-07 peta0 = 9.831615184e-14
+ etab = -5.692749632e-01 letab = 1.007241565e-07 wetab = 4.799240839e-07 petab = -8.920348947e-14
+ u0 = 6.180697291e-02 lu0 = -1.066579166e-08 wu0 = -5.081970886e-08 pu0 = 9.445859286e-15
+ ua = 3.236330670e-09 lua = -9.377386158e-16 wua = -4.468080755e-15 pua = 8.304821699e-22
+ ub = 1.960605889e-18 lub = -2.214160605e-26 wub = -1.054997168e-25 pub = 1.960923236e-32
+ uc = 2.470670693e-12 luc = -4.432691369e-19 wuc = -2.112056181e-18 puc = 3.925678823e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.162674144e+06 lvsat = 2.267196024e-01 wvsat = 1.080259597e+00 pvsat = -2.007878512e-7
+ a0 = 8.484088001e+00 la0 = -1.366290969e-06 wa0 = -6.510019672e-06 pa0 = 1.210017356e-12
+ ags = 1.249999978e+00 lags = 5.733106434e-15 wags = 6.674690667e-14 pags = -1.240625380e-20
+ a1 = 0.0
+ a2 = -4.887798307e+00 la2 = 1.028419613e-06 wa2 = 4.900150830e-06 pa2 = -9.107910348e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.480033014e-02 lketa = -8.183149155e-09 wketa = -3.899045977e-08 pketa = 7.247156758e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.169231343e-01 lpclm = 9.579261270e-10 wpclm = 4.564207222e-09 ppclm = -8.483491964e-16
+ pdiblc1 = 6.690069315e-01 lpdiblc1 = -9.317227188e-08 wpdiblc1 = -4.439416121e-07 ppdiblc1 = 8.251542744e-14
+ pdiblc2 = 3.900619837e-02 lpdiblc2 = -6.532799657e-09 wpdiblc2 = -3.112709477e-08 ppdiblc2 = 5.785593105e-15
+ pdiblcb = -1.826808881e+00 lpdiblcb = 2.689764300e-07 wpdiblcb = 1.281601909e-06 ppdiblcb = -2.382113468e-13
+ drout = 1.000002240e+00 ldrout = -3.873937047e-13 wdrout = -1.128322708e-12 pdrout = 2.097213425e-19
+ pscbe1 = 8.000000120e+08 lpscbe1 = -2.218666077e-06 wpscbe1 = -1.030905151e-05 ppscbe1 = 1.916145325e-12
+ pscbe2 = -2.553424115e-08 lpscbe2 = 6.117437060e-15 wpscbe2 = 2.914798799e-14 ppscbe2 = -5.417736528e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.253625129e+01 lbeta0 = -7.778277127e-07 wbeta0 = -3.706147693e-06 pbeta0 = 6.888616717e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.428176633e-08 lagidl = -1.004673247e-14 wagidl = -4.787005594e-14 pagidl = 8.897607298e-21
+ bgidl = 1.000000279e+09 lbgidl = -4.367739868e-05 wbgidl = -7.342895508e-06 pbgidl = 1.364822388e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 4.927942511e-01 lkt1 = -1.912721729e-07 wkt1 = -9.113619559e-07 pkt1 = 1.693948467e-13
+ kt2 = -9.625899344e-02 lkt2 = -1.726053078e-15 wkt2 = -2.076593475e-14 pkt2 = 3.859764064e-21
+ at = 6.929996725e+05 lat = -1.211390386e-01 wat = -5.771958716e-01 pat = 1.072833967e-7
+ ute = -1.593596795e+00 lute = 2.869083286e-07 wute = 1.367043055e-06 pute = -2.540922926e-13
+ ua1 = 7.435796928e-10 lua1 = 3.355629547e-23 wua1 = -4.230078833e-22 pua1 = 7.862447675e-29
+ ub1 = -4.726027072e-19 lub1 = 4.829925600e-31 wub1 = 1.801473603e-30 pub1 = -3.348398998e-37
+ uc1 = -2.193903712e-11 luc1 = 6.556618174e-24 wuc1 = 2.276894790e-23 puc1 = -4.232064257e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.108 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.109 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.110389418e+00 lvth0 = 3.885659956e-7
+ k1 = 4.210956021e-01 lk1 = 2.110826255e-7
+ k2 = 1.775005695e-02 lk2 = 2.994270855e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 3.388131789e-27 pcit = 3.794707604e-31
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.944604484e-01 lvoff = 4.898018407e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.149046479e+00 lnfactor = -5.147691351e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.179692641e-02 lu0 = -1.779462005e-8
+ ua = -8.962599665e-10 lua = 1.912151425e-15 wua = 6.617444900e-30
+ ub = 1.670762721e-18 lub = -5.162101108e-24
+ uc = -1.282222813e-10 luc = 4.509347416e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.679434283e+04 lvsat = 1.066639228e+0
+ a0 = 1.543433334e+00 la0 = -1.587782595e-6
+ ags = 8.823956664e-02 lags = 5.007298559e-7
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-06 wa2 = 7.105427358e-21
+ b0 = -1.712879585e-07 lb0 = 1.368397233e-12
+ b1 = 3.860850241e-09 lb1 = -3.084383066e-14
+ keta = 4.015882949e-02 lketa = -3.357644528e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 wpclm = 1.110223025e-22 ppclm = -6.217248938e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.914844237e-03 lpdiblc2 = -1.274661131e-8
+ pdiblcb = -2.715221659e-01 lpdiblcb = 9.299255256e-7
+ drout = 0.56
+ pscbe1 = 8.000324548e+08 lpscbe1 = -6.487344658e-1
+ pscbe2 = 1.314643402e-08 lpscbe2 = -6.168183535e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.579227219e+01 lbeta0 = -3.156696758e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.869014186e-09 lagidl = -1.936435346e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.229045954e-01 legidl = 1.045227198e-05 wegidl = 8.881784197e-22 pegidl = -2.131628207e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365713387e-01 lkt1 = -3.355454267e-08 wkt1 = -3.552713679e-21
+ kt2 = -6.266527973e-02 lkt2 = 8.233974711e-8
+ at = 1.182508234e+05 lat = -9.446904559e-1
+ ute = -5.016829954e-02 lute = -6.558688149e-7
+ ua1 = 2.268269050e-09 lua1 = -3.559399084e-15
+ ub1 = -1.570431596e-18 lub1 = 6.826830664e-24
+ uc1 = -4.378798232e-11 luc1 = 2.798238376e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.110 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-1
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595753e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 ppdiblc2 = -2.775557562e-29
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+3
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 wpscbe2 = -5.293955920e-29
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.111 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569065e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077654e-03 lketa = -3.715224604e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = -1.332267630e-21 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048848e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807946e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123884e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.112 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-08 pk2 = -2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-06 pdsub = 3.552713679e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = -2.775557562e-22 peta0 = 3.469446952e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = -5.412337245e-22 petab = 2.116362641e-27
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-9
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16 pagidl = 1.654361225e-36
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = -3.552713679e-21 pute = 5.329070518e-27
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.113 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.060692995e+00 lvth0 = 2.691011409e-8
+ k1 = 5.224851534e-01 lk1 = -6.227372655e-9
+ k2 = -7.144540537e-03 lk2 = 3.224478319e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.223655613e+00 ldsub = -4.419034005e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.288458330e-01 lvoff = 1.026340558e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.087125419e+00 lnfactor = -4.927330750e-7
+ eta0 = -7.462418332e-03 leta0 = 2.249307616e-7
+ etab = -1.632744345e+00 letab = 7.978799692e-7
+ u0 = 1.148561965e-02 lu0 = -2.566038196e-9
+ ua = -1.059609635e-10 lua = -5.351404061e-16
+ ub = 4.864006036e-19 lub = 3.665394455e-25
+ uc = -9.754060033e-11 luc = 3.244585840e-17 wuc = -8.271806126e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.249860650e+04 lvsat = 3.449316359e-2
+ a0 = 1.648107076e+00 la0 = -4.403606970e-7
+ ags = -3.625107541e-01 lags = 7.883081323e-7
+ a1 = 0.0
+ a2 = 1.047418086e+00 la2 = -4.690021102e-8
+ b0 = -8.575503616e-17 lb0 = 8.480058261e-23
+ b1 = -3.565229431e-20 lb1 = 3.525548427e-26
+ keta = 1.023393023e-02 lketa = -2.366260124e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.536347840e+00 lpclm = -7.221227228e-7
+ pdiblc1 = 6.191336573e-02 lpdiblc1 = -2.265833997e-8
+ pdiblc2 = 7.533057929e-04 lpdiblc2 = -3.197073994e-10
+ pdiblcb = -1.477237207e-02 lpdiblcb = -1.011379443e-8
+ drout = 1.036997061e+00 ldrout = -3.658528362e-8
+ pscbe1 = 8.230739141e+08 lpscbe1 = -3.636238561e+1
+ pscbe2 = 3.809477986e-09 lpscbe2 = 5.307539814e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.632459620e+00 lbeta0 = 1.024241563e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.004804533e-09 lagidl = -4.912187918e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.254810687e-01 lkt1 = -5.298728500e-8
+ kt2 = -6.206186670e-02 lkt2 = 1.335240081e-8
+ at = 8.443425409e+04 lat = -2.242016604e-2
+ ute = -1.875821105e+00 lute = 8.184494349e-7
+ ua1 = -3.292299871e-09 lua1 = 2.830042980e-15 wua1 = -6.617444900e-30
+ ub1 = 4.034982618e-18 lub1 = -3.105147788e-24 pub1 = 6.162975822e-45
+ uc1 = 3.136276955e-10 luc1 = -2.439630433e-16 wuc1 = -8.271806126e-31 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.114 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.809317576e-01 lvth0 = -1.208276190e-8
+ k1 = 4.446623754e-01 lk1 = 3.181784882e-8
+ k2 = 1.132757422e-02 lk2 = -5.805984424e-09 wk2 = -2.081668171e-23 pk2 = -1.214306433e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.244403898e-01 ldsub = 2.171402925e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.700309796e-01 lvoff = -1.848941181e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.825934693e-01 lnfactor = 5.361094594e-7
+ eta0 = 4.169452362e-01 leta0 = 1.745059157e-8
+ etab = -1.210426333e-03 letab = 2.719825911e-10
+ u0 = 4.591262030e-03 lu0 = 8.044064145e-10
+ ua = -1.330850367e-09 lua = 6.367127645e-17
+ ub = 7.875179014e-19 lub = 2.193322321e-25
+ uc = -6.000952568e-11 luc = 1.409804193e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.833766079e+04 lvsat = -2.582274881e-3
+ a0 = 8.732071908e-01 la0 = -6.153539006e-8
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 1.100021230e+00 la2 = -7.261631000e-8
+ b0 = 1.715100723e-16 lb0 = -4.096861098e-23
+ b1 = 7.130458861e-20 lb1 = -1.703252708e-26
+ keta = -4.438001254e-02 lketa = 3.036516966e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.930264200e-01 lpclm = 2.699774716e-07 wpclm = -1.776356839e-21 ppclm = -8.881784197e-28
+ pdiblc1 = -3.561786926e-01 lpdiblc1 = 1.817343246e-07 wpdiblc1 = -6.661338148e-22 ppdiblc1 = 3.330669074e-28
+ pdiblc2 = -8.000440691e-03 lpdiblc2 = 3.959736644e-09 wpdiblc2 = -2.428612866e-23 ppdiblc2 = -1.062518129e-29
+ pdiblcb = 2.058549522e-01 lpdiblcb = -1.179718745e-07 ppdiblcb = -4.440892099e-28
+ drout = 1.376341573e+00 ldrout = -2.024806355e-7
+ pscbe1 = 6.996965507e+08 lpscbe1 = 2.395310605e+1
+ pscbe2 = 2.022856548e-08 lpscbe2 = -2.719259489e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.553332902e+00 lbeta0 = 8.518424213e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.492459760e-12 lagidl = 7.296188029e-19
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.443546811e-01 lkt1 = 5.126457872e-9
+ kt2 = -1.748919269e-02 lkt2 = -8.437842332e-9
+ at = 1.056349506e+04 lat = 1.369303193e-2
+ ute = 4.030997005e-01 lute = -2.956465794e-07 pute = 8.881784197e-28
+ ua1 = 4.600244176e-09 lua1 = -1.028385029e-15
+ ub1 = -4.368480081e-18 lub1 = 1.003053022e-24
+ uc1 = -2.690313562e-10 luc1 = 4.088148730e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.115 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 1.892511455e+00 lvth0 = -6.984621420e-07 wvth0 = -2.378273038e-06 pvth0 = 5.680980805e-13
+ k1 = -1.023469066e+00 lk1 = 3.825104063e-07 wk1 = 2.797392848e-07 pk1 = -6.682132296e-14
+ k2 = -1.230143196e+00 lk2 = 2.907441384e-07 wk2 = 1.515881498e-06 pk2 = -3.620986135e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.935836715e+00 ldsub = -5.138680996e-07 wdsub = -8.906975653e-07 pdsub = 2.127609274e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.856935526e-01 lvoff = 9.138907021e-09 wvoff = 2.755572190e-07 pvoff = -6.582235290e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 4.639453174e+00 lnfactor = -3.374046181e-07 wnfactor = -2.146745620e-06 pnfactor = 5.127931263e-13
+ eta0 = 3.379817246e+00 leta0 = -6.902906454e-07 weta0 = -1.981322228e-06 peta0 = 4.732784405e-13
+ etab = 2.804513364e-01 letab = -6.700856268e-08 wetab = -1.901181056e-07 petab = 4.541351189e-14
+ u0 = 6.253850934e-03 lu0 = 4.072638031e-10 wu0 = 9.062285602e-09 pu0 = -2.164708162e-15
+ ua = -1.075622216e-09 lua = 2.704928080e-18 wua = 1.600658304e-15 pua = -3.823492491e-22
+ ub = 3.218834943e-18 lub = -3.614364695e-25 wub = -1.630086402e-24 pub = 3.893787388e-31
+ uc = -1.122147664e-10 luc = 2.656830778e-17 wuc = 9.620518080e-17 puc = -2.298053154e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.602221845e+05 lvsat = -4.364033106e-02 wvsat = -1.181578322e-01 pvsat = 2.822436138e-8
+ a0 = -2.751867379e+00 la0 = 8.043861723e-07 wa0 = 1.876227659e-06 pa0 = -4.481745008e-13
+ ags = 2.122259388e+00 lags = -1.472984433e-07 wags = -2.419574230e-14 pags = 5.779632772e-21
+ a1 = 0.0
+ a2 = 1.997655719e+00 la2 = -2.870342606e-07 wa2 = -7.419762549e-07 pa2 = 1.772358680e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.201734676e-01 lketa = 4.502829959e-08 wketa = 9.763195825e-08 pketa = -2.332134587e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.631235178e-01 lpclm = -6.192064035e-09 wpclm = 9.355739020e-09 ppclm = -2.234805380e-15
+ pdiblc1 = 2.492799844e+00 lpdiblc1 = -4.988011784e-07 wpdiblc1 = -1.343193772e-06 ppdiblc1 = 3.208486964e-13
+ pdiblc2 = -1.269330109e-03 lpdiblc2 = 2.351876259e-09 wpdiblc2 = 1.879854120e-08 ppdiblc2 = -4.490407537e-15
+ pdiblcb = -6.214551482e+00 lpdiblcb = 1.415670610e-06 wpdiblcb = 5.444514951e-06 ppdiblcb = -1.300531286e-12
+ drout = -6.083433780e-01 ldrout = 2.716010589e-07 wdrout = 1.091991919e-12 pdrout = -2.608441108e-19
+ pscbe1 = 7.999088766e+08 lpscbe1 = 1.538776180e-02 wpscbe1 = -3.270675659e-06 ppscbe1 = 7.812652588e-13
+ pscbe2 = -5.619405608e-09 lpscbe2 = 3.455045365e-15 wpscbe2 = 1.594294487e-14 ppscbe2 = -3.808291240e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.027741067e+01 lbeta0 = -3.266462140e-07 wbeta0 = -1.784425886e-08 pbeta0 = 4.262458114e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.434877663e-08 lagidl = 5.816565390e-15 wagidl = 2.107863972e-14 pagidl = -5.035054671e-21
+ bgidl = 1.818113554e+09 lbgidl = -1.381548295e+02 wbgidl = -1.213946533e-05 pbgidl = 2.899753571e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.076005616e-01 lkt1 = 9.189500134e-08 wkt1 = 3.692842564e-07 pkt1 = -8.821093032e-14
+ kt2 = 4.201323668e-01 lkt2 = -1.129725043e-07 wkt2 = -3.260290076e-07 pkt2 = 7.787854904e-14
+ at = -5.390357964e+04 lat = 2.909228206e-02 wat = 1.647532354e-01 pat = -3.935460534e-8
+ ute = -6.234815451e+00 lute = 1.289952213e-06 wute = 3.106286707e-06 pute = -7.419987058e-13
+ ua1 = -3.973509631e-09 lua1 = 1.019627543e-15 wua1 = 2.822004629e-15 pua1 = -6.740922457e-22
+ ub1 = 3.466488140e-18 lub1 = -8.684858370e-25 wub1 = -2.571998166e-24 pub1 = 6.143732019e-31
+ uc1 = -3.407032927e-10 luc1 = 5.800176276e-17 wuc1 = 5.278353894e-17 puc1 = -1.260840395e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.116 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -6.706882806e+00 lvth0 = 8.295936765e-07 wvth0 = 4.938638984e-06 pvth0 = -7.347064039e-13
+ k1 = 1.241650052e+00 lk1 = -2.851902678e-13 wk1 = -1.159590357e-07 pk1 = 2.778285619e-19
+ k2 = 2.953107055e+00 lk2 = -4.575276194e-07 wk2 = -2.808362802e-06 pk2 = 4.051965135e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.071503902e-01 ldsub = 1.246905478e-12 wdsub = 3.692163642e-07 pdsub = -8.121330382e-19
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.315756283e-01 lvoff = 1.445490305e-14 wvoff = -1.142239185e-07 pvoff = -1.343579115e-20
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.641432990e+00 lnfactor = 1.156073893e-12 wnfactor = 8.898732738e-07 pnfactor = -7.774339679e-19
+ eta0 = -7.078861471e-01 leta0 = -1.908779499e-13 weta0 = 8.212970885e-07 peta0 = 1.283245954e-19
+ etab = -1.163551493e-01 letab = 1.635138200e-13 wetab = 7.880833243e-08 petab = -1.053403134e-19
+ u0 = -2.382875480e-02 lu0 = 6.039716633e-09 wu0 = 2.502117559e-08 pu0 = -5.348906382e-15
+ ua = -1.059671604e-09 lua = 1.249060394e-20 wua = -6.634466295e-16 pua = -1.084047267e-26
+ ub = 1.078507955e-18 lub = 6.041441199e-31 wub = 6.757056197e-25 pub = -3.961149418e-37
+ uc = 4.511518326e-11 luc = -9.001619704e-25 wuc = -3.987897469e-17 puc = -2.200399853e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.694732941e+05 lvsat = -6.834007000e-02 wvsat = -2.766438816e-01 pvsat = 6.052348596e-8
+ a0 = 2.011474541e+00 la0 = 6.849440410e-13 wa0 = -7.777307944e-07 pa0 = -5.909088330e-19
+ ags = 1.249999985e+00 lags = 2.209453953e-15 wags = 5.998725783e-14 pags = -9.285635372e-21
+ a1 = 0.0
+ a2 = 2.979207143e-01 la2 = -1.129221872e-14 wa2 = 3.075639787e-07 pa2 = 9.650872101e-21
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.647176683e-02 lketa = -8.932938632e-14 wketa = -4.047072088e-08 pketa = 5.894958298e-20
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.264555378e-01 lpclm = 6.356443194e-14 wpclm = -3.877899051e-09 ppclm = -4.503795026e-20
+ pdiblc1 = -4.609599909e-01 lpdiblc1 = 2.695344090e-13 wpdiblc1 = 5.567819536e-07 ppdiblc1 = -2.250310684e-19
+ pdiblc2 = 1.265778096e-02 lpdiblc2 = 5.518142804e-15 wpdiblc2 = -7.792356648e-09 ppdiblc2 = -2.880564148e-21
+ pdiblcb = 2.168643790e+00 lpdiblcb = 4.676120611e-13 wpdiblcb = -2.256858877e-06 ppdiblcb = -3.170625238e-19
+ drout = 1.000004036e+00 ldrout = -6.261631498e-13 wdrout = -2.718649313e-12 pdrout = 4.211808147e-19
+ pscbe1 = 7.999999866e+08 lpscbe1 = 2.216106415e-06 wpscbe1 = 1.217721558e-05 ppscbe1 = -2.011379242e-12
+ pscbe2 = 1.484038863e-08 lpscbe2 = -9.757385448e-23 wpscbe2 = -6.608672385e-15 ppscbe2 = 4.017563031e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.343098775e+00 lbeta0 = 1.139656035e-12 wbeta0 = 7.400419436e-09 pbeta0 = -6.721896284e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.009526615e-08 lagidl = -1.271299343e-22 wagidl = -8.737519279e-15 pagidl = 1.100464676e-28
+ bgidl = 1.000000297e+09 lbgidl = -4.814885712e-05 wbgidl = -2.361618042e-05 pbgidl = 5.324844360e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.634238901e-01 lkt1 = -1.245555694e-13 wkt1 = -1.530763332e-07 pkt1 = 1.127552736e-19
+ kt2 = -2.488580142e-01 lkt2 = -1.085374475e-13 wkt2 = 1.351450292e-07 pkt2 = 9.845428472e-20
+ at = 1.183725023e+05 lat = 2.212370769e-08 wat = -6.829340789e-02 pat = -2.056943020e-14
+ ute = 1.403913598e+00 lute = 4.218140015e-14 wute = -1.287618094e-06 pute = -2.156912648e-21
+ ua1 = 2.064428120e-09 lua1 = 1.095570711e-21 wua1 = -1.169772848e-15 pua1 = -8.619188631e-28
+ ub1 = -1.676437835e-18 lub1 = 7.956157116e-32 wub1 = 1.066144675e-24 pub1 = 2.244745922e-38
+ uc1 = 2.766521061e-12 luc1 = 1.686011016e-23 wuc1 = -2.187976307e-17 puc1 = -1.335706324e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.117 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.118 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.110389418e+00 lvth0 = 3.885659956e-7
+ k1 = 4.210956021e-01 lk1 = 2.110826255e-7
+ k2 = 1.775005695e-02 lk2 = 2.994270855e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 pcit = -1.897353802e-31
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.944604484e-01 lvoff = 4.898018407e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.149046479e+00 lnfactor = -5.147691352e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.179692641e-02 lu0 = -1.779462005e-8
+ ua = -8.962599665e-10 lua = 1.912151425e-15
+ ub = 1.670762721e-18 lub = -5.162101108e-24
+ uc = -1.282222813e-10 luc = 4.509347416e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.679434283e+04 lvsat = 1.066639228e+0
+ a0 = 1.543433334e+00 la0 = -1.587782595e-6
+ ags = 8.823956664e-02 lags = 5.007298559e-7
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = -1.712879585e-07 lb0 = 1.368397233e-12
+ b1 = 3.860850241e-09 lb1 = -3.084383066e-14
+ keta = 4.015882949e-02 lketa = -3.357644528e-07 pketa = 8.881784197e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.914844237e-03 lpdiblc2 = -1.274661131e-8
+ pdiblcb = -2.715221659e-01 lpdiblcb = 9.299255256e-7
+ drout = 0.56
+ pscbe1 = 8.000324548e+08 lpscbe1 = -6.487344658e-1
+ pscbe2 = 1.314643402e-08 lpscbe2 = -6.168183535e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.579227219e+01 lbeta0 = -3.156696758e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.869014186e-09 lagidl = -1.936435346e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.229045954e-01 legidl = 1.045227198e-05 pegidl = -7.105427358e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365713387e-01 lkt1 = -3.355454267e-8
+ kt2 = -6.266527973e-02 lkt2 = 8.233974711e-8
+ at = 1.182508234e+05 lat = -9.446904559e-1
+ ute = -5.016829954e-02 lute = -6.558688149e-7
+ ua1 = 2.268269050e-09 lua1 = -3.559399084e-15
+ ub1 = -1.570431596e-18 lub1 = 6.826830664e-24
+ uc1 = -4.378798232e-11 luc1 = 2.798238376e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.119 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-01 pvsat = -3.725290298e-21
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595752e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-08 wpdiblc2 = -1.734723476e-24 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+3
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17 wuc1 = -5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.120 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569066e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077653e-03 lketa = -3.715224604e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = 8.881784197e-22 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048849e-01 lkt1 = 2.502969993e-8
+ kt2 = -6.021807946e-02 lkt2 = 1.562472077e-8
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123884e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.121 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-06 pdsub = 1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = -3.434752482e-22 peta0 = -1.838806885e-28
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = 1.543903894e-21 petab = 3.268219029e-27
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-9
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16 pagidl = -8.271806126e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = -8.881784197e-22 pute = -1.332267630e-27
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24 pub1 = -1.232595164e-44
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.122 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.060692995e+00 lvth0 = 2.691011409e-8
+ k1 = 5.224851534e-01 lk1 = -6.227372655e-9
+ k2 = -7.144540537e-03 lk2 = 3.224478319e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.223655613e+00 ldsub = -4.419034005e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.288458330e-01 lvoff = 1.026340558e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.087125419e+00 lnfactor = -4.927330750e-07 wnfactor = -1.421085472e-20
+ eta0 = -7.462418332e-03 leta0 = 2.249307616e-7
+ etab = -1.632744345e+00 letab = 7.978799692e-7
+ u0 = 1.148561965e-02 lu0 = -2.566038196e-9
+ ua = -1.059609635e-10 lua = -5.351404061e-16
+ ub = 4.864006036e-19 lub = 3.665394455e-25
+ uc = -9.754060033e-11 luc = 3.244585840e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.249860650e+04 lvsat = 3.449316359e-2
+ a0 = 1.648107076e+00 la0 = -4.403606970e-7
+ ags = -3.625107541e-01 lags = 7.883081323e-07 pags = 1.776356839e-27
+ a1 = 0.0
+ a2 = 1.047418086e+00 la2 = -4.690021102e-8
+ b0 = -8.575503616e-17 lb0 = 8.480058261e-23
+ b1 = -3.565229431e-20 lb1 = 3.525548427e-26
+ keta = 1.023393023e-02 lketa = -2.366260124e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.536347840e+00 lpclm = -7.221227228e-7
+ pdiblc1 = 6.191336573e-02 lpdiblc1 = -2.265833997e-8
+ pdiblc2 = 7.533057929e-04 lpdiblc2 = -3.197073994e-10
+ pdiblcb = -1.477237207e-02 lpdiblcb = -1.011379443e-8
+ drout = 1.036997061e+00 ldrout = -3.658528362e-8
+ pscbe1 = 8.230739141e+08 lpscbe1 = -3.636238561e+1
+ pscbe2 = 3.809477986e-09 lpscbe2 = 5.307539814e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.632459620e+00 lbeta0 = 1.024241563e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.004804533e-09 lagidl = -4.912187918e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.254810687e-01 lkt1 = -5.298728500e-8
+ kt2 = -6.206186670e-02 lkt2 = 1.335240081e-8
+ at = 8.443425409e+04 lat = -2.242016604e-2
+ ute = -1.875821105e+00 lute = 8.184494349e-7
+ ua1 = -3.292299871e-09 lua1 = 2.830042980e-15 wua1 = 3.308722450e-30 pua1 = 3.308722450e-36
+ ub1 = 4.034982618e-18 lub1 = -3.105147788e-24 wub1 = 6.162975822e-39
+ uc1 = 3.136276955e-10 luc1 = -2.439630433e-16 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.123 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.809317576e-01 lvth0 = -1.208276190e-8
+ k1 = 4.446623754e-01 lk1 = 3.181784882e-8
+ k2 = 1.132757422e-02 lk2 = -5.805984424e-09 wk2 = -2.081668171e-23 pk2 = -9.540979118e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.244403898e-01 ldsub = 2.171402925e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.700309796e-01 lvoff = -1.848941181e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.825934693e-01 lnfactor = 5.361094594e-7
+ eta0 = 4.169452362e-01 leta0 = 1.745059157e-8
+ etab = -1.210426333e-03 letab = 2.719825911e-10
+ u0 = 4.591262030e-03 lu0 = 8.044064145e-10
+ ua = -1.330850367e-09 lua = 6.367127645e-17 wua = -6.617444900e-30
+ ub = 7.875179014e-19 lub = 2.193322321e-25
+ uc = -6.000952568e-11 luc = 1.409804193e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.833766079e+04 lvsat = -2.582274881e-3
+ a0 = 8.732071908e-01 la0 = -6.153539006e-8
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 1.100021230e+00 la2 = -7.261631000e-8
+ b0 = 1.715100723e-16 lb0 = -4.096861098e-23
+ b1 = 7.130458861e-20 lb1 = -1.703252708e-26
+ keta = -4.438001254e-02 lketa = 3.036516966e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.930264200e-01 lpclm = 2.699774716e-07 wpclm = -4.440892099e-22 ppclm = 4.440892099e-28
+ pdiblc1 = -3.561786926e-01 lpdiblc1 = 1.817343246e-07 wpdiblc1 = -6.661338148e-22 ppdiblc1 = -1.942890293e-28
+ pdiblc2 = -8.000440691e-03 lpdiblc2 = 3.959736644e-09 ppdiblc2 = -5.204170428e-30
+ pdiblcb = 2.058549522e-01 lpdiblcb = -1.179718745e-7
+ drout = 1.376341573e+00 ldrout = -2.024806355e-07 wdrout = -7.105427358e-21
+ pscbe1 = 6.996965507e+08 lpscbe1 = 2.395310605e+1
+ pscbe2 = 2.022856548e-08 lpscbe2 = -2.719259489e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.553332902e+00 lbeta0 = 8.518424213e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.492459760e-12 lagidl = 7.296188029e-19
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.443546811e-01 lkt1 = 5.126457872e-9
+ kt2 = -1.748919269e-02 lkt2 = -8.437842332e-9
+ at = 1.056349506e+04 lat = 1.369303193e-2
+ ute = 4.030997005e-01 lute = -2.956465794e-07 pute = 4.440892099e-28
+ ua1 = 4.600244176e-09 lua1 = -1.028385029e-15 wua1 = 1.323488980e-29
+ ub1 = -4.368480081e-18 lub1 = 1.003053022e-24
+ uc1 = -2.690313562e-10 luc1 = 4.088148730e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.124 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.549615042e-01 lvth0 = -4.217327634e-8
+ k1 = -7.003034297e-01 lk1 = 3.053158307e-7
+ k2 = 5.210617164e-01 lk2 = -1.275661790e-07 pk2 = 1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.906868453e+00 ldsub = -2.680784508e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.264079998e-02 lvoff = -6.690161979e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.159449638e+00 lnfactor = 2.549938263e-7
+ eta0 = 1.090917209e+00 leta0 = -1.435410936e-7
+ etab = 6.081955074e-02 letab = -1.454511803e-08 wetab = -8.500145032e-23 petab = 1.669671346e-29
+ u0 = 1.672295362e-02 lu0 = -2.093490755e-9
+ ua = 7.735201398e-10 lua = -4.389997064e-16
+ ub = 1.335696111e-18 lub = 8.838890319e-26
+ uc = -1.074822148e-12 luc = 2.030929986e-20
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.237216887e+05 lvsat = -1.103445762e-2
+ a0 = -5.843766510e-01 la0 = 2.866376622e-7
+ ags = 2.122259360e+00 lags = -1.472984366e-7
+ a1 = 0.0
+ a2 = 1.140496064e+00 la2 = -8.228453375e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.073852549e-01 lketa = 1.808657922e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.739316293e-01 lpclm = -8.773797609e-9
+ pdiblc1 = 9.410904691e-01 lpdiblc1 = -1.281443601e-7
+ pdiblc2 = 2.044747146e-02 lpdiblc2 = -2.835616130e-9
+ pdiblcb = 7.516267856e-02 lpdiblcb = -8.675341105e-8
+ drout = -6.083421165e-01 ldrout = 2.716007575e-7
+ pscbe1 = 7.999088728e+08 lpscbe1 = 1.538866434e-2
+ pscbe2 = 1.279850067e-08 lpscbe2 = -9.444399071e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025679629e+01 lbeta0 = -3.217220576e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.082891577e-12 lagidl = -1.244253710e-19
+ bgidl = 1.818113540e+09 lbgidl = -1.381548261e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.809891118e-01 lkt1 = -1.000967566e-8
+ kt2 = 4.349105275e-02 lkt2 = -2.300419356e-8
+ at = 1.364257274e+05 lat = -1.637167951e-2
+ ute = -2.646312955e+00 lute = 4.327666216e-7
+ ua1 = -7.134207826e-10 lua1 = 2.408901201e-16
+ ub1 = 4.952164236e-19 lub1 = -1.587381621e-25
+ uc1 = -2.797257078e-10 luc1 = 4.343604708e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.125 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.244846545e-01 lvth0 = -7.067055642e-08 wvth0 = -2.398564691e-07 pvth0 = 4.458212191e-14
+ k1 = 4.084085152e-01 lk1 = 1.299754278e-07 wk1 = 6.053131695e-07 pk1 = -1.125095588e-13
+ k2 = -3.370385465e-01 lk2 = 1.908693761e-08 wk2 = 3.965961450e-08 pk2 = -7.371532548e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.545913526e+00 ldsub = -4.138449893e-07 wdsub = -1.927334129e-06 pdsub = 3.582335946e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.049129247e+00 lvoff = 1.274320494e-07 wvoff = 5.934684802e-07 pvoff = -1.103079864e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.010648547e+00 lnfactor = -9.927685021e-07 wnfactor = -4.623459835e-06 pnfactor = 8.593624796e-13
+ eta0 = 5.170531424e+00 leta0 = -9.162691482e-07 weta0 = -4.267190487e-06 peta0 = 7.931426957e-13
+ etab = 4.499375087e-01 letab = -8.833471760e-08 wetab = -4.113870507e-07 petab = 7.646451112e-14
+ u0 = -3.699187191e-03 lu0 = 1.491622615e-09 wu0 = 7.596579014e-09 pu0 = -1.411976141e-15
+ ua = -5.808584233e-09 lua = 7.402223043e-16 wua = 3.447316618e-15 pua = -6.407527398e-22
+ ub = 5.914965134e-18 lub = -7.538617939e-25 wub = -3.510838116e-24 pub = 6.525594806e-31
+ uc = -2.414450447e-10 luc = 4.469996709e-17 wuc = 2.081738630e-16 puc = -3.869327591e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.754167315e+05 lvsat = 4.345557102e-02 wvsat = 1.950249121e-01 pvsat = -3.624928042e-8
+ a0 = -3.555136077e+00 la0 = 8.676682875e-07 wa0 = 4.040849822e-06 pa0 = -7.510727564e-13
+ ags = 1.250000055e+00 lags = -8.517666572e-15
+ a1 = 0.0
+ a2 = 2.507997991e+00 la2 = -3.447456312e-07 wa2 = -1.605527534e-06 pa2 = 2.984194027e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.431940821e-01 lketa = 4.515012654e-08 wketa = 2.102704106e-07 pketa = -3.908296121e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.985881834e-01 lpclm = 4.347037898e-09 wpclm = 2.024469605e-08 ppclm = -3.762881655e-15
+ pdiblc1 = 3.539925496e+00 lpdiblc1 = -6.240900108e-07 wpdiblc1 = -2.906472543e-06 ppdiblc1 = 5.402260516e-13
+ pdiblc2 = -4.333623387e-02 lpdiblc2 = 8.734402102e-09 wpdiblc2 = 4.067729445e-08 ppdiblc2 = -7.560688720e-15
+ pdiblcb = -1.404858519e+01 lpdiblcb = 2.529694214e-06 wpdiblcb = 1.178113131e-05 ppdiblcb = -2.189758877e-12
+ drout = 1.000000895e+00 ldrout = -1.395987859e-13
+ pscbe1 = 8.000000007e+08 lpscbe1 = -1.075172424e-7
+ pscbe2 = -3.264784285e-08 lpscbe2 = 7.407595996e-15 wpscbe2 = 3.449818553e-14 ppscbe2 = -6.412177744e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.396250352e+00 lbeta0 = -8.289871313e-09 wbeta0 = -3.860875508e-08 pbeta0 = 7.176209307e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.433070876e-10 lagidl = -4.497329248e-17 wagidl = -2.094467713e-16 pagidl = 3.892987138e-23
+ bgidl = 1.000000270e+09 lbgidl = -4.199738693e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.459058749e+00 lkt1 = 1.707764623e-07 wkt1 = 7.953293048e-07 pkt1 = -1.478278579e-13
+ kt2 = 7.222637721e-01 lkt2 = -1.514834916e-07 wkt2 = -7.054793537e-07 pkt2 = 1.311274475e-13
+ at = -3.723674392e+05 lat = 7.654958324e-02 wat = 3.565018818e-01 pat = -6.626300477e-8
+ ute = -7.848584152e+00 lute = 1.443279018e-06 wute = 6.721547513e-06 pute = -1.249334036e-12
+ ua1 = -6.341296857e-09 lua1 = 1.311193651e-15 wua1 = 6.106407618e-15 pua1 = -1.134997984e-21
+ ub1 = 5.984608789e-18 lub1 = -1.195031558e-24 wub1 = -5.565425826e-24 pub1 = 1.034445698e-30
+ uc1 = -1.544564348e-10 luc1 = 2.452491740e-17 wuc1 = 1.142158864e-16 puc1 = -2.122930681e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.126 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.127 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.110389418e+00 lvth0 = 3.885659956e-07 wvth0 = -3.552713679e-21
+ k1 = 4.210956021e-01 lk1 = 2.110826255e-7
+ k2 = 1.775005695e-02 lk2 = 2.994270855e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 5.082197684e-27 pcit = -2.710505431e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.944604484e-01 lvoff = 4.898018407e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.149046479e+00 lnfactor = -5.147691352e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.179692641e-02 lu0 = -1.779462005e-8
+ ua = -8.962599665e-10 lua = 1.912151425e-15
+ ub = 1.670762721e-18 lub = -5.162101108e-24
+ uc = -1.282222813e-10 luc = 4.509347416e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.679434284e+04 lvsat = 1.066639228e+0
+ a0 = 1.543433334e+00 la0 = -1.587782595e-6
+ ags = 8.823956664e-02 lags = 5.007298559e-7
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = -1.712879585e-07 lb0 = 1.368397233e-12
+ b1 = 3.860850240e-09 lb1 = -3.084383066e-14
+ keta = 4.015882949e-02 lketa = -3.357644528e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.914844237e-03 lpdiblc2 = -1.274661131e-8
+ pdiblcb = -2.715221659e-01 lpdiblcb = 9.299255256e-7
+ drout = 0.56
+ pscbe1 = 8.000324548e+08 lpscbe1 = -6.487344657e-1
+ pscbe2 = 1.314643402e-08 lpscbe2 = -6.168183535e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.579227219e+01 lbeta0 = -3.156696758e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.869014186e-09 lagidl = -1.936435346e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.229045954e-01 legidl = 1.045227198e-05 pegidl = -7.105427358e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365713387e-01 lkt1 = -3.355454267e-8
+ kt2 = -6.266527973e-02 lkt2 = 8.233974711e-8
+ at = 1.182508234e+05 lat = -9.446904559e-1
+ ute = -5.016829954e-02 lute = -6.558688149e-7
+ ua1 = 2.268269050e-09 lua1 = -3.559399084e-15
+ ub1 = -1.570431596e-18 lub1 = 6.826830664e-24
+ uc1 = -4.378798232e-11 luc1 = 2.798238376e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.128 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.067909815e+00 lvth0 = 4.920197463e-8
+ k1 = 4.556026508e-01 lk1 = -6.458970099e-8
+ k2 = 1.888114602e-02 lk2 = 2.090658503e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.249456820e-01 lvoff = -6.554259092e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.646126736e+00 lnfactor = -4.022586465e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.241315721e-03 lu0 = 2.621821543e-9
+ ua = -6.951832022e-10 lua = 3.057752950e-16
+ ub = 1.032606613e-18 lub = -6.395491904e-26
+ uc = -7.084610619e-11 luc = -7.436062681e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.668846287e+05 lvsat = -8.514108537e-1
+ a0 = 1.377626083e+00 la0 = -2.631700178e-7
+ ags = 8.902569586e-02 lags = 4.944495718e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.453595753e-04 lketa = -8.187316924e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398542052e-01 lpclm = -7.900610979e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.382883923e-03 lpdiblc2 = 1.359851026e-8
+ pdiblcb = -2.485894473e-01 lpdiblcb = 7.467190179e-7
+ drout = 0.56
+ pscbe1 = 1.223533045e+09 lpscbe1 = -3.383939895e+3
+ pscbe2 = -1.692187543e-08 lpscbe2 = 1.785299800e-13 wpscbe2 = -2.646977960e-29
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.454111638e+00 lbeta0 = 2.256438486e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.898162607e-10 lagidl = -1.955024528e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.668713786e+00 legidl = -6.257395361e-06 pegidl = -1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.064088808e-01 lkt1 = -2.745184978e-7
+ kt2 = -4.842691408e-02 lkt2 = -3.140870509e-8
+ at = -9.042369403e+04 lat = 7.223831365e-1
+ ute = -1.644424595e-01 lute = 2.570525935e-7
+ ua1 = 5.811130231e-10 lua1 = 9.919071081e-15
+ ub1 = 8.106627581e-19 lub1 = -1.219542258e-23 pub1 = -1.232595164e-44
+ uc1 = -1.162365659e-11 luc1 = 2.286722078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.129 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058035232e+00 lvth0 = 9.813546376e-9
+ k1 = 4.427490850e-01 lk1 = -1.331849770e-8
+ k2 = 2.173134058e-02 lk2 = 9.537529476e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.570387389e-01 ldsub = -1.184848914e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.653962750e-01 lvoff = 9.580956600e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 8.357297946e-01 lnfactor = 3.198851581e-6
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391144744e-01 letab = 2.756886533e-7
+ u0 = 8.885569066e-03 lu0 = 4.040848704e-9
+ ua = -7.590571481e-10 lua = 5.605601617e-16
+ ub = 1.009458227e-18 lub = 2.838098239e-26
+ uc = -7.555427377e-11 luc = 1.134420574e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.332582857e+00 la0 = -8.349844430e-8
+ ags = 1.492824772e-01 lags = 2.540931044e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.416077653e-03 lketa = -3.715224604e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.457365877e-01 lpclm = 2.343558448e-06 wpclm = -6.661338148e-22 ppclm = -2.220446049e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.613575983e-03 lpdiblc2 = -6.331718765e-9
+ pdiblcb = -9.757511029e-02 lpdiblcb = 1.443424596e-7
+ drout = 0.56
+ pscbe1 = -3.954447050e+07 lpscbe1 = 1.654312115e+3
+ pscbe2 = 4.621586901e-08 lpscbe2 = -7.331827470e-14 wpscbe2 = 1.058791184e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.143313392e+01 lbeta0 = -9.262897737e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.687073149e-10 lagidl = -2.752756878e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815048848e-01 lkt1 = 2.502969993e-08 wkt1 = 1.776356839e-21
+ kt2 = -6.021807947e-02 lkt2 = 1.562472077e-08 wkt2 = 2.220446049e-22
+ at = 1.020960915e+05 lat = -4.555326054e-2
+ ute = -1.321769333e-01 lute = 1.283496039e-7
+ ua1 = 3.319292612e-09 lua1 = -1.003171333e-15
+ ub1 = -2.832123884e-18 lub1 = 2.335179770e-24
+ uc1 = 1.777277470e-11 luc1 = -9.439132211e-17 wuc1 = -2.584939414e-32 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.130 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.072503618e+00 lvth0 = 3.858928540e-8
+ k1 = 3.568093539e-01 lk1 = 1.576044552e-7
+ k2 = 5.659888429e-02 lk2 = -5.980948219e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.484432034e-01 ldsub = 1.013810956e-06 pdsub = 1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.159937502e-01 lvoff = -2.445633576e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.300976860e+00 lnfactor = 2.846656514e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = 1.734723476e-22 peta0 = -7.979727989e-29
+ etab = 8.156999796e-01 letab = -1.623313170e-06 wetab = 5.655198532e-22 petab = 1.307981501e-27
+ u0 = 1.292134394e-02 lu0 = -3.985782875e-9
+ ua = -3.091838044e-10 lua = -3.341794354e-16
+ ub = 1.188535755e-18 lub = -3.277809421e-25
+ uc = -7.491430767e-11 luc = 1.007139638e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.942857446e+04 lvsat = -1.191447383e-2
+ a0 = 1.377432675e+00 la0 = -1.726989017e-7
+ ags = 1.211644219e-01 lags = 3.100162610e-7
+ a1 = 0.0
+ a2 = 6.022358887e-01 la2 = 3.933271080e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.084892703e-02 lketa = -2.814396178e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.610337555e-01 lpclm = 3.412231158e-7
+ pdiblc1 = 7.370933700e-01 lpdiblc1 = -6.903235908e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.248972000e-01 ldrout = 8.653629058e-7
+ pscbe1 = 7.981125877e+08 lpscbe1 = -1.167887878e+1
+ pscbe2 = 9.524462383e-09 lpscbe2 = -3.438368068e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.893237408e+00 lbeta0 = 1.755236233e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.432540367e-10 lagidl = 7.429488855e-16 pagidl = 8.271806126e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.588881710e-01 lkt1 = -1.995200383e-8
+ kt2 = -5.612249362e-02 lkt2 = 7.479132955e-9
+ at = 9.642825824e+04 lat = -3.428067692e-2
+ ute = 9.019606480e-01 lute = -1.928415607e-06 wute = -8.881784197e-22 pute = 4.440892099e-28
+ ua1 = 6.024083757e-09 lua1 = -6.382649298e-15
+ ub1 = -4.182471934e-18 lub1 = 5.020846495e-24 pub1 = 6.162975822e-45
+ uc1 = -1.252175596e-10 luc1 = 1.899978642e-16 wuc1 = 2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.131 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.060692995e+00 lvth0 = 2.691011409e-8
+ k1 = 5.224851534e-01 lk1 = -6.227372655e-9
+ k2 = -7.144540537e-03 lk2 = 3.224478319e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.223655613e+00 ldsub = -4.419034005e-07 wdsub = -3.552713679e-21
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.288458330e-01 lvoff = 1.026340558e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.087125419e+00 lnfactor = -4.927330750e-7
+ eta0 = -7.462418332e-03 leta0 = 2.249307616e-7
+ etab = -1.632744345e+00 letab = 7.978799692e-7
+ u0 = 1.148561965e-02 lu0 = -2.566038196e-9
+ ua = -1.059609635e-10 lua = -5.351404061e-16
+ ub = 4.864006036e-19 lub = 3.665394455e-25
+ uc = -9.754060033e-11 luc = 3.244585840e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.249860650e+04 lvsat = 3.449316359e-2
+ a0 = 1.648107076e+00 la0 = -4.403606970e-7
+ ags = -3.625107541e-01 lags = 7.883081323e-07 pags = -8.881784197e-28
+ a1 = 0.0
+ a2 = 1.047418086e+00 la2 = -4.690021102e-8
+ b0 = -8.575503616e-17 lb0 = 8.480058261e-23
+ b1 = -3.565229431e-20 lb1 = 3.525548427e-26
+ keta = 1.023393023e-02 lketa = -2.366260124e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.536347840e+00 lpclm = -7.221227228e-7
+ pdiblc1 = 6.191336573e-02 lpdiblc1 = -2.265833997e-8
+ pdiblc2 = 7.533057929e-04 lpdiblc2 = -3.197073994e-10
+ pdiblcb = -1.477237207e-02 lpdiblcb = -1.011379443e-8
+ drout = 1.036997061e+00 ldrout = -3.658528362e-8
+ pscbe1 = 8.230739141e+08 lpscbe1 = -3.636238561e+1
+ pscbe2 = 3.809477986e-09 lpscbe2 = 5.307539814e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.632459620e+00 lbeta0 = 1.024241563e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.004804533e-09 lagidl = -4.912187918e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.254810687e-01 lkt1 = -5.298728500e-8
+ kt2 = -6.206186670e-02 lkt2 = 1.335240081e-08 wkt2 = -2.220446049e-22
+ at = 8.443425409e+04 lat = -2.242016604e-2
+ ute = -1.875821105e+00 lute = 8.184494349e-7
+ ua1 = -3.292299871e-09 lua1 = 2.830042980e-15 wua1 = -3.308722450e-30 pua1 = -1.654361225e-36
+ ub1 = 4.034982618e-18 lub1 = -3.105147788e-24 pub1 = -3.081487911e-45
+ uc1 = 3.136276955e-10 luc1 = -2.439630433e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.132 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.809317576e-01 lvth0 = -1.208276190e-8
+ k1 = 4.446623754e-01 lk1 = 3.181784882e-8
+ k2 = 1.132757422e-02 lk2 = -5.805984424e-09 wk2 = 3.469446952e-24 pk2 = -6.071532166e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.244403898e-01 ldsub = 2.171402925e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.700309796e-01 lvoff = -1.848941181e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.825934693e-01 lnfactor = 5.361094594e-7
+ eta0 = 4.169452362e-01 leta0 = 1.745059157e-8
+ etab = -1.210426333e-03 letab = 2.719825911e-10
+ u0 = 4.591262030e-03 lu0 = 8.044064145e-10
+ ua = -1.330850367e-09 lua = 6.367127645e-17
+ ub = 7.875179014e-19 lub = 2.193322321e-25
+ uc = -6.000952568e-11 luc = 1.409804193e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.833766079e+04 lvsat = -2.582274881e-3
+ a0 = 8.732071908e-01 la0 = -6.153539006e-8
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 1.100021230e+00 la2 = -7.261631000e-8
+ b0 = 1.715100723e-16 lb0 = -4.096861098e-23
+ b1 = 7.130458861e-20 lb1 = -1.703252708e-26
+ keta = -4.438001254e-02 lketa = 3.036516966e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.930264200e-01 lpclm = 2.699774716e-07 ppclm = -3.330669074e-28
+ pdiblc1 = -3.561786926e-01 lpdiblc1 = 1.817343246e-07 wpdiblc1 = -3.330669074e-22 ppdiblc1 = 1.387778781e-29
+ pdiblc2 = -8.000440691e-03 lpdiblc2 = 3.959736644e-09 wpdiblc2 = -4.336808690e-25 ppdiblc2 = 6.830473687e-30
+ pdiblcb = 2.058549522e-01 lpdiblcb = -1.179718745e-07 ppdiblcb = 5.551115123e-29
+ drout = 1.376341573e+00 ldrout = -2.024806355e-7
+ pscbe1 = 6.996965507e+08 lpscbe1 = 2.395310605e+1
+ pscbe2 = 2.022856548e-08 lpscbe2 = -2.719259489e-15 wpscbe2 = -5.293955920e-29
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.553332902e+00 lbeta0 = 8.518424213e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.492459760e-12 lagidl = 7.296188029e-19
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.443546811e-01 lkt1 = 5.126457872e-9
+ kt2 = -1.748919269e-02 lkt2 = -8.437842332e-9
+ at = 1.056349506e+04 lat = 1.369303193e-2
+ ute = 4.030997005e-01 lute = -2.956465794e-7
+ ua1 = 4.600244176e-09 lua1 = -1.028385029e-15
+ ub1 = -4.368480081e-18 lub1 = 1.003053022e-24
+ uc1 = -2.690313562e-10 luc1 = 4.088148730e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.133 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.549615042e-01 lvth0 = -4.217327634e-8
+ k1 = -7.003034297e-01 lk1 = 3.053158307e-7
+ k2 = 5.210617164e-01 lk2 = -1.275661790e-07 wk2 = 4.440892099e-22 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.906868453e+00 ldsub = -2.680784508e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.264079998e-02 lvoff = -6.690161979e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.159449638e+00 lnfactor = 2.549938263e-7
+ eta0 = 1.090917209e+00 leta0 = -1.435410936e-07 weta0 = 3.552713679e-21
+ etab = 6.081955074e-02 letab = -1.454511803e-08 wetab = -5.898059818e-23 petab = -1.138412281e-29
+ u0 = 1.672295362e-02 lu0 = -2.093490755e-9
+ ua = 7.735201398e-10 lua = -4.389997064e-16
+ ub = 1.335696111e-18 lub = 8.838890319e-26
+ uc = -1.074822148e-12 luc = 2.030929986e-20
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.237216887e+05 lvsat = -1.103445762e-2
+ a0 = -5.843766510e-01 la0 = 2.866376622e-7
+ ags = 2.122259360e+00 lags = -1.472984366e-7
+ a1 = 0.0
+ a2 = 1.140496064e+00 la2 = -8.228453375e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.073852549e-01 lketa = 1.808657922e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.739316293e-01 lpclm = -8.773797609e-9
+ pdiblc1 = 9.410904691e-01 lpdiblc1 = -1.281443601e-7
+ pdiblc2 = 2.044747146e-02 lpdiblc2 = -2.835616130e-9
+ pdiblcb = 7.516267856e-02 lpdiblcb = -8.675341105e-8
+ drout = -6.083421165e-01 ldrout = 2.716007575e-7
+ pscbe1 = 7.999088728e+08 lpscbe1 = 1.538866434e-2
+ pscbe2 = 1.279850067e-08 lpscbe2 = -9.444399071e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025679629e+01 lbeta0 = -3.217220576e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.082891577e-12 lagidl = -1.244253710e-19
+ bgidl = 1.818113540e+09 lbgidl = -1.381548261e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.809891118e-01 lkt1 = -1.000967566e-8
+ kt2 = 4.349105275e-02 lkt2 = -2.300419356e-8
+ at = 1.364257274e+05 lat = -1.637167951e-2
+ ute = -2.646312955e+00 lute = 4.327666216e-7
+ ua1 = -7.134207826e-10 lua1 = 2.408901201e-16 pua1 = 4.135903063e-37
+ ub1 = 4.952164236e-19 lub1 = -1.587381621e-25 pub1 = -1.925929944e-46
+ uc1 = -2.797257078e-10 luc1 = 4.343604708e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.134 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -7.751851307e-01 lvth0 = -6.124685891e-08 wvth0 = -1.974900358e-07 pvth0 = 3.670747295e-14
+ k1 = 4.032537413e-01 lk1 = 1.309335456e-07 wk1 = 6.096206119e-07 pk1 = -1.133101831e-13
+ k2 = -1.270326679e-01 lk2 = -1.994685504e-08 wk2 = -1.358259178e-07 pk2 = 2.524596334e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.562326471e+00 ldsub = -4.168956634e-07 wdsub = -1.941049147e-06 pdsub = 3.607828049e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.049131121e+00 lvoff = 1.274323978e-07 wvoff = 5.934700462e-07 pvoff = -1.103082775e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.010648022e+00 lnfactor = -9.927684046e-07 wnfactor = -4.623459397e-06 pnfactor = 8.593623981e-13
+ eta0 = 5.170532605e+00 leta0 = -9.162693676e-07 weta0 = -4.267191473e-06 peta0 = 7.931428791e-13
+ etab = 4.534408311e-01 letab = -8.898588015e-08 wetab = -4.143145040e-07 petab = 7.700863687e-14
+ u0 = -2.271727163e-03 lu0 = 1.226300619e-09 wu0 = 6.403762010e-09 pu0 = -1.190267245e-15
+ ua = -5.808672994e-09 lua = 7.402388024e-16 wua = 3.447390789e-15 pua = -6.407665260e-22
+ ub = 5.914943214e-18 lub = -7.538577197e-25 wub = -3.510819799e-24 pub = 6.525560761e-31
+ uc = -2.432178282e-10 luc = 4.502947436e-17 wuc = 2.096552399e-16 puc = -3.896861943e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.916160934e+04 lvsat = 2.184723147e-02 wvsat = 9.787957447e-02 pvsat = -1.819287651e-8
+ a0 = -3.555135937e+00 la0 = 8.676682617e-07 wa0 = 4.040849706e-06 pa0 = -7.510727348e-13
+ ags = 1.250000055e+00 lags = -8.517666572e-15
+ a1 = 0.0
+ a2 = 2.521670470e+00 la2 = -3.472869348e-07 wa2 = -1.616952558e-06 pa2 = 3.005429719e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.431940735e-01 lketa = 4.515012496e-08 wketa = 2.102704034e-07 pketa = -3.908295989e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.984157820e-01 lpclm = 4.379082144e-09 wpclm = 2.038875844e-08 ppclm = -3.789658532e-15
+ pdiblc1 = 3.564676665e+00 lpdiblc1 = -6.286905107e-07 wpdiblc1 = -2.927155165e-06 ppdiblc1 = 5.440703305e-13
+ pdiblc2 = -4.368263680e-02 lpdiblc2 = 8.798788014e-09 wpdiblc2 = 4.096675636e-08 ppdiblc2 = -7.614491005e-15
+ pdiblcb = -1.414891189e+01 lpdiblcb = 2.548341936e-06 wpdiblcb = 1.186496650e-05 ppdiblcb = -2.205341324e-12
+ drout = 1.000000895e+00 ldrout = -1.395988072e-13 wdrout = -8.526512829e-20 pdrout = 1.421085472e-26
+ pscbe1 = 8.000000007e+08 lpscbe1 = -1.075172424e-7
+ pscbe2 = -3.294162523e-08 lpscbe2 = 7.462201327e-15 wpscbe2 = 3.474367655e-14 ppscbe2 = -6.457807160e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.396579140e+00 lbeta0 = -8.350983044e-09 wbeta0 = -3.888349715e-08 pbeta0 = 7.227275615e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.368158513e-10 lagidl = -2.517976639e-17 wagidl = -1.204603515e-16 pagidl = 2.238996552e-23
+ bgidl = 1.000000270e+09 lbgidl = -4.199739456e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.459059860e+00 lkt1 = 1.707766687e-07 wkt1 = 7.953302329e-07 pkt1 = -1.478280304e-13
+ kt2 = 7.282715491e-01 lkt2 = -1.526001571e-07 wkt2 = -7.104995844e-07 pkt2 = 1.320605577e-13
+ at = -3.754033662e+05 lat = 7.711387099e-02 wat = 3.590387691e-01 pat = -6.673453602e-8
+ ute = -7.905824039e+00 lute = 1.453918196e-06 wute = 6.769378422e-06 pute = -1.258224367e-12
+ ua1 = -6.393298287e-09 lua1 = 1.320859156e-15 wua1 = 6.149861156e-15 pua1 = -1.143074693e-21
+ ub1 = 6.032003283e-18 lub1 = -1.203840772e-24 wub1 = -5.605029708e-24 pub1 = 1.041806872e-30
+ uc1 = -1.554290835e-10 luc1 = 2.470570361e-17 wuc1 = 1.150286531e-16 puc1 = -2.138037575e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.135 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.136 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.136723888e+00 lvth0 = 9.149622934e-07 wvth0 = 2.095228371e-08 pvth0 = -4.188124752e-13
+ k1 = 4.806021126e-01 lk1 = -9.783852781e-07 wk1 = -4.734468894e-08 pk1 = 9.463668324e-13
+ k2 = -3.958080703e-02 lk2 = 1.175921896e-06 wk2 = 4.561369666e-08 pk2 = -9.117662528e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 8.470329473e-28 pcit = -8.131516294e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -4.993651811e-01 lvoff = 4.585615905e-06 wvoff = 1.630267133e-07 pvoff = -3.258719778e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.641082999e+00 lnfactor = 7.570892850e-05 wnfactor = 3.015510395e-06 pnfactor = -6.027664528e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.629416808e-02 lu0 = -1.076893991e-07 wu0 = -3.578104410e-09 pu0 = 7.152226390e-14
+ ua = -7.744305291e-10 lua = -5.230813610e-16 wua = -9.693018063e-17 pua = 1.937524780e-21
+ ub = 1.229356260e-18 lub = 3.661115263e-24 wub = 3.511926915e-25 pub = -7.019945055e-30
+ uc = -4.796256430e-10 luc = 7.475090855e-15 wuc = 2.795842454e-16 puc = -5.588573135e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.584995976e+05 lvsat = 2.076155172e+01 wvsat = 7.839215355e-01 pvsat = -1.566970566e-5
+ a0 = 3.147366166e-01 la0 = 2.297247637e-05 wa0 = 9.775781400e-07 pa0 = -1.954068236e-11
+ ags = -2.772122112e-01 lags = 7.805697935e-06 wags = 2.907614744e-07 pags = -5.811993313e-12
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = 5.968156421e-07 lb0 = -1.398512579e-11 wb0 = -6.111201230e-13 pb0 = 1.221560069e-17
+ b1 = 1.083324021e-08 lb1 = -1.702140274e-13 wb1 = -5.547386855e-15 pb1 = 1.108859947e-19
+ keta = 1.295143122e-01 lketa = -2.121879580e-06 wketa = -7.109318784e-08 pketa = 1.421072490e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 ppclm = 1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.033233594e-03 lpdiblc2 = -1.511308078e-08 wpdiblc2 = -9.419317700e-11 ppdiblc2 = 1.882815170e-15
+ pdiblcb = -9.652811730e-01 lpdiblcb = 1.479738413e-05 wpdiblcb = 5.519699288e-07 ppdiblcb = -1.103325515e-11
+ drout = 0.56
+ pscbe1 = 8.005164348e+08 lpscbe1 = -1.032294826e+01 wpscbe1 = -3.850651552e-01 ppscbe1 = 7.697017329e-6
+ pscbe2 = 7.697886426e-08 lpscbe2 = -1.337619985e-12 wpscbe2 = -5.078648581e-14 ppscbe2 = 1.015164463e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 1.324310849e+01 lbeta0 = 3.349513260e-04 wbeta0 = 2.589683072e-05 pbeta0 = -5.176483827e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.778694999e-09 lagidl = -3.754784497e-14 wagidl = -7.237620677e-16 pagidl = 1.446718588e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -8.220688001e+00 legidl = 1.663211508e-04 wegidl = 6.204088029e-06 pegidl = -1.240127091e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.203490209e-01 lkt1 = -2.356707345e-06 wkt1 = -9.246903295e-08 pkt1 = 1.848351479e-12
+ kt2 = -2.494669610e-02 lkt2 = -6.716121177e-07 wkt2 = -3.000973495e-08 pkt2 = 5.998606906e-13
+ at = 7.314087702e+05 lat = -1.320102494e+01 wat = -4.878419519e-01 pat = 9.751409357e-6
+ ute = -9.142973343e+00 lute = 1.810990291e-04 wute = 7.234435734e-06 pute = -1.446081954e-10
+ ua1 = -2.010032758e-08 lua1 = 4.435635709e-13 wua1 = 1.779694758e-14 pua1 = -3.557408716e-19
+ ub1 = 1.442100735e-17 lub1 = -3.128239635e-22 wub1 = -1.272314063e-23 pub1 = 2.543212041e-28
+ uc1 = 7.075481051e-10 luc1 = -1.473853554e-14 wuc1 = -5.977795205e-16 puc1 = 1.194893712e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.137 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.054859051e+00 lvth0 = 2.609547583e-07 wvth0 = -1.038347492e-08 pvth0 = -1.684751732e-13
+ k1 = 3.847944230e-01 lk1 = -2.129901005e-07 wk1 = 5.633658385e-08 pk1 = 1.180706227e-13
+ k2 = 7.103734872e-02 lk2 = 2.922078298e-07 wk2 = -4.149662230e-08 pk2 = -2.158532389e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 4.212900146e-01 lvoff = -2.769378767e-06 wvoff = -5.141593374e-07 pvoff = 2.151231546e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.522810662e+01 lnfactor = -1.389455344e-04 wnfactor = -1.796672000e-05 pnfactor = 1.073476656e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.560547132e-02 lu0 = -1.021874902e-07 wu0 = -5.063462207e-09 pu0 = 8.338859424e-14
+ ua = 1.585742728e-09 lua = -1.937819869e-14 wua = -1.814754850e-15 pua = 1.566100275e-20
+ ub = 6.987221940e-19 lub = 7.900281830e-24 wub = 2.656457888e-25 pub = -6.336521971e-30
+ uc = 4.684238456e-10 luc = -9.875326261e-17 wuc = -4.290550376e-16 puc = 7.265397324e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.301030589e+06 lvsat = -1.326728120e+01 wvsat = -2.414033277e+00 pvsat = 9.878339601e-6
+ a0 = 4.479082834e+00 la0 = -1.029594420e-05 wa0 = -2.467587223e-06 pa0 = 7.982295860e-12
+ ags = 7.401130783e-01 lags = -3.215815508e-07 wags = -5.180194454e-07 pags = 6.492523138e-13
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -8.932513360e-07 lb0 = -2.081174407e-12 wb0 = 7.106904144e-13 pb0 = 1.655828144e-18
+ b1 = 1.348973816e-08 lb1 = -1.914364441e-13 wb1 = -1.073273245e-14 pb1 = 1.523110466e-19
+ keta = -1.258448413e-01 lketa = -8.184849989e-08 wketa = 9.945233762e-08 pketa = 5.860645772e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.873812691e+00 lpclm = -7.775450302e-05 wpclm = -7.664989318e-06 ppclm = 6.123460321e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -2.547549491e-02 lpdiblc2 = 2.046505751e-07 wpdiblc2 = 1.916861134e-08 ppdiblc2 = -1.520052259e-13
+ pdiblcb = -6.003656642e-01 lpdiblcb = 1.188212157e-05 wpdiblcb = 2.798808973e-07 ppdiblcb = -8.859571249e-12
+ drout = 0.56
+ pscbe1 = 7.539444167e+09 lpscbe1 = -5.384674054e+04 wpscbe1 = -5.025077838e+03 ppscbe1 = 4.014931437e-2
+ pscbe2 = -4.871533919e-07 lpscbe2 = 3.169159272e-12 wpscbe2 = 3.741265396e-13 ppscbe2 = -2.379410459e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.387094614e-09 lalpha0 = 1.188020555e-14 walpha0 = 1.183165191e-15 palpha0 = -9.452152897e-21
+ alpha1 = -1.387094614e-09 lalpha1 = 1.188020555e-14 walpha1 = 1.183165191e-15 palpha1 = -9.452152897e-21
+ beta0 = 4.117415699e+02 lbeta0 = -2.848601077e-03 wbeta0 = -3.248424841e-04 pbeta0 = 2.284362407e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.382417225e-10 lagidl = -1.245917200e-14 wagidl = 4.103383728e-17 pagidl = 8.357330821e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 2.506206400e+01 legidl = -9.957042824e-05 wegidl = -1.861226409e-05 pegidl = 7.424190184e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.943739230e-01 lkt1 = -2.564219025e-06 wkt1 = -8.913747720e-08 pkt1 = 1.821736113e-12
+ kt2 = -1.949679391e-01 lkt2 = 6.866654895e-07 wkt2 = 1.165912634e-07 pkt2 = -5.713156268e-13
+ at = -1.776518596e+06 lat = 6.834480753e+00 wat = 1.341494198e+00 pat = -4.862919330e-6
+ ute = 2.587998156e+01 lute = -9.869480461e-05 wute = -2.072151673e-05 pute = 7.872827453e-11
+ ua1 = 5.314906596e-08 lua1 = -1.416163116e-13 wua1 = -4.182421985e-14 pua1 = 1.205648842e-19
+ ub1 = -3.054091048e-17 lub1 = 4.637095299e-23 wub1 = 2.494400140e-23 pub1 = -4.659669686e-29
+ uc1 = -8.396166079e-09 luc1 = 5.798985360e-14 wuc1 = 6.670926411e-15 puc1 = -4.611980963e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.138 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.767428606e-01 lvth0 = -5.064057157e-08 wvth0 = -6.467799929e-08 pvth0 = 4.809862623e-14
+ k1 = 1.283183924e+00 lk1 = -3.796549029e-06 wk1 = -6.686684474e-07 pk1 = 3.010021442e-12
+ k2 = -2.143982826e-01 lk2 = 1.430773456e-06 wk2 = 1.878699230e-07 pk2 = -1.130766571e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.377755770e-01 ldsub = -1.108010666e-06 wdsub = 1.532619541e-08 pdsub = -6.113420107e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -5.220727687e-01 lvoff = 9.935727378e-07 wvoff = 2.042174653e-07 pvoff = -7.142801303e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.959945825e+01 lnfactor = 3.986579434e-05 wnfactor = 1.625868519e-05 pnfactor = -2.917302633e-11
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391329935e-01 letab = 2.757625239e-07 wetab = 1.473425771e-11 petab = -5.877303857e-17
+ u0 = -2.708917017e-02 lu0 = 6.811588438e-08 wu0 = 2.862229398e-08 pu0 = -5.097950803e-14
+ ua = -6.190868297e-09 lua = 1.164169173e-14 wua = 4.321668450e-15 pua = -8.816392061e-21
+ ub = 2.570623141e-18 lub = 4.335123017e-25 wub = -1.242097151e-24 pub = -3.223313906e-31
+ uc = 7.864042300e-10 luc = -1.367135679e-15 wuc = -6.857931487e-16 puc = 1.096748923e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.942369141e+05 lvsat = 1.472660479e+00 wvsat = 3.561800105e-01 pvsat = -1.171681076e-6
+ a0 = 3.486131913e-01 la0 = 6.179962244e-06 wa0 = 7.828679131e-07 pa0 = -4.983347120e-12
+ ags = 2.978324380e+00 lags = -9.249515467e-06 wags = -2.250847977e-06 pags = 7.561280059e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.125184709e-06 lb0 = -1.156022336e-12 wb0 = 8.952217082e-13 pb0 = 9.197568027e-19
+ b1 = -9.297840862e-08 lb1 = 2.332511525e-13 wb1 = 7.397566743e-14 pb1 = -1.855797485e-19
+ keta = -2.339630630e-01 lketa = 3.494210314e-07 wketa = 1.912509327e-07 pketa = -3.075662042e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.774215065e+01 lpclm = 3.240198468e-05 wpclm = 1.368184535e-05 ppclm = -2.391514520e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 5.125638564e-02 lpdiblc2 = -1.014229212e-07 wpdiblc2 = -3.790566750e-08 ppdiblc2 = 7.565665270e-14
+ pdiblcb = 4.768531366e+00 lpdiblcb = -9.533710729e-06 wpdiblcb = -3.871581367e-06 ppdiblcb = 7.700072034e-12
+ drout = 0.56
+ pscbe1 = -1.255920101e+10 lpscbe1 = 2.632414227e+04 wpscbe1 = 9.960914179e+03 ppscbe1 = -1.962785960e-2
+ pscbe2 = 6.053861159e-07 lpscbe2 = -1.188838794e-12 wpscbe2 = -4.448881502e-13 ppscbe2 = 8.875326668e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.074189227e-09 lalpha0 = -5.915275728e-15 walpha0 = -2.366330381e-15 palpha0 = 4.706323505e-21
+ alpha1 = 3.074189227e-09 lalpha1 = -5.915275728e-15 walpha1 = -2.366330381e-15 palpha1 = 4.706323505e-21
+ beta0 = -6.277588731e+02 lbeta0 = 1.297831055e-03 wbeta0 = 5.085552230e-04 pbeta0 = -1.039952705e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.256001918e-09 lagidl = -3.087881711e-14 wagidl = -3.968001307e-15 pagidl = 2.434885084e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.164895998e+00 lkt1 = 9.081803661e-07 wkt1 = 5.437210046e-07 pkt1 = -7.026540994e-13
+ kt2 = -1.677425974e-02 lkt2 = -2.412593213e-08 wkt2 = -3.456485874e-08 pkt2 = 3.162649396e-14
+ at = -7.852348418e+05 lat = 2.880378726e+00 wat = 7.059800118e-01 pat = -2.327935859e-6
+ ute = -7.147168510e-01 lute = 7.387990047e-06 wute = 4.634815744e-07 pute = -5.775929648e-12
+ ua1 = 9.969868771e-09 lua1 = 3.061989271e-14 wua1 = -5.291344705e-15 pua1 = -2.516000546e-20
+ ub1 = -1.685864092e-17 lub1 = -8.205841577e-24 wub1 = 1.115980554e-23 pub1 = 8.386668487e-30
+ uc1 = 1.324591417e-08 luc1 = -2.833759103e-14 wuc1 = -1.052460031e-14 puc1 = 2.247091104e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.139 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.454862106e-01 lvth0 = -1.128059850e-07 wvth0 = -1.010578439e-07 pvth0 = 1.204534078e-13
+ k1 = -1.875322662e+00 lk1 = 2.485309964e-06 wk1 = 1.775933339e-06 pk1 = -1.851973712e-12
+ k2 = 9.789291513e-01 lk2 = -9.425996770e-07 wk2 = -7.338262517e-07 pk2 = 7.023673004e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -7.830572264e+00 ldsub = 1.613220630e-05 wdsub = 6.032508687e-06 pdsub = -1.202852794e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.090911116e-01 lvoff = 1.722059096e-07 wvoff = -8.505409107e-08 pvoff = -1.389566100e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.419813634e-01 lnfactor = -5.906846742e-07 wnfactor = 1.240371115e-06 pnfactor = 6.964479767e-13
+ eta0 = 3.764988462e+00 leta0 = -7.487078167e-06 weta0 = -3.167805135e-06 peta0 = 6.300352600e-12
+ etab = 1.297621799e+01 letab = -2.580896558e-05 wetab = -9.675175659e-06 petab = 1.924263714e-11
+ u0 = 1.509192283e-02 lu0 = -1.577682605e-08 wu0 = -1.726960315e-09 pu0 = 9.381213353e-15
+ ua = -7.635836457e-10 lua = 8.475281065e-16 wua = 3.615305106e-16 pua = -9.401925179e-22
+ ub = 6.477219506e-18 lub = -7.336200012e-24 wub = -4.207793143e-24 pub = 5.576052397e-30
+ uc = 5.727359548e-10 luc = -9.421772562e-16 wuc = -5.152847972e-16 puc = 7.576299775e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.070857726e+05 lvsat = -7.177271727e-01 wvsat = -5.152903153e-01 pvsat = 5.615601111e-7
+ a0 = 6.486720840e+00 la0 = -6.027935915e-06 wa0 = -4.065062068e-06 pa0 = 4.658555383e-12
+ ags = -1.844703121e+00 lags = 3.428592389e-07 wags = 1.564087466e-06 pags = -2.613059573e-14
+ a1 = 0.0
+ a2 = -2.346909555e+00 la2 = 6.258794007e-06 wa2 = 2.346404996e-06 pa2 = -4.666694505e-12
+ b0 = -1.821158003e-06 lb0 = 2.281780713e-13 wb0 = 1.448953373e-12 pb0 = -1.815434934e-19
+ b1 = 1.876228144e-07 lb1 = -3.248282019e-13 wb1 = -1.492768388e-13 pb1 = 2.584404636e-19
+ keta = 8.430415854e-02 lketa = -2.835710976e-07 wketa = -7.570588825e-08 pketa = 2.233762083e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.307511939e+00 lpclm = 9.659974780e-06 wpclm = 5.385203862e-06 ppclm = -7.414203836e-12
+ pdiblc1 = 5.829624753e+00 lpdiblc1 = -1.081870648e-05 wpdiblc1 = -4.051730004e-06 ppdiblc1 = 8.058364253e-12
+ pdiblc2 = 9.415235240e-05 lpdiblc2 = 3.321096633e-10 wpdiblc2 = 2.672077771e-10 ppdiblc2 = -2.642337545e-16
+ pdiblcb = -2.974292909e+00 lpdiblcb = 5.865760187e-06 wpdiblcb = 2.346522322e-06 ppdiblcb = -4.666927852e-12
+ drout = -3.762780049e+00 ldrout = 8.597447556e-06 wdrout = 3.093121548e-06 pdrout = -6.151816653e-12
+ pscbe1 = 7.699666654e+08 lpscbe1 = -1.858394578e+02 wpscbe1 = 2.239351502e+01 ppscbe1 = 1.385659882e-4
+ pscbe2 = 6.023023057e-09 lpscbe2 = 3.216480191e-15 wpscbe2 = 2.785822160e-15 ppscbe2 = -2.832666530e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.406692809e+01 lbeta0 = 1.434273567e-06 wbeta0 = -1.445938813e-05 pbeta0 = 2.553649582e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.022105960e-08 lagidl = -9.695377140e-17 wagidl = 7.938561618e-15 pagidl = 6.682450317e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.349135889e-01 lkt1 = 4.507752512e-07 wkt1 = 3.787362950e-07 pkt1 = -3.745209601e-13
+ kt2 = -9.469036779e-03 lkt2 = -3.865507092e-08 wkt2 = -3.711851664e-08 pkt2 = 3.670538755e-14
+ at = 1.110109726e+06 lat = -8.892152242e-01 wat = -8.065072765e-01 pat = 6.802047344e-7
+ ute = 7.003004925e+00 lute = -7.961555261e-06 wute = -4.854125050e-06 pute = 4.800098638e-12
+ ua1 = 5.087427921e-08 lua1 = -5.073366207e-14 wua1 = -3.568380220e-14 pua1 = 3.528664149e-20
+ ub1 = -4.321027080e-17 lub1 = 4.420412454e-23 wub1 = 3.105137539e-23 pub1 = -3.117507805e-29
+ uc1 = -2.059363702e-09 luc1 = 2.102616960e-15 wuc1 = 1.538849222e-15 puc1 = -1.521721830e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.140 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.112276128e+00 lvth0 = 5.212756031e-08 wvth0 = 4.104067542e-08 pvth0 = -2.006355499e-14
+ k1 = 7.633193985e-01 lk1 = -1.239640101e-07 wk1 = -1.916130238e-07 pk1 = 9.367385893e-14
+ k2 = 5.140453207e-02 lk2 = -2.539840681e-08 wk2 = -4.658293025e-08 pk2 = 2.277299711e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.646496638e+01 ldsub = -7.892922996e-06 wdsub = -1.212632216e-05 pdsub = 5.928195113e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.318828776e-01 lvoff = -2.638600392e-07 wvoff = -4.461280982e-07 pvoff = 2.180986434e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.746862984e+00 lnfactor = 1.870458836e-06 wnfactor = 3.846027522e-06 pnfactor = -1.880207475e-12
+ eta0 = -7.970553271e+00 leta0 = 4.117846987e-06 weta0 = 6.335610271e-06 peta0 = -3.097289793e-12
+ etab = -2.595370628e+01 letab = 1.268766863e-05 wetab = 1.935029238e-05 petab = -9.459777436e-12
+ u0 = -7.803626012e-03 lu0 = 6.863895332e-09 wu0 = 1.534694821e-08 pu0 = -7.502662573e-15
+ ua = 1.358769378e-09 lua = -1.251203128e-15 wua = -1.165371684e-15 pua = 5.697152551e-22
+ ub = -3.070796135e-18 lub = 2.105546215e-24 wub = 2.830183984e-24 pub = -1.383592044e-30
+ uc = -7.211540753e-10 luc = 3.373117779e-16 wuc = 4.961606002e-16 puc = -2.425580326e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.182292441e+05 lvsat = 9.840208790e-02 wvsat = 1.040099539e-01 pvsat = -5.084734617e-8
+ a0 = 4.247662510e-02 la0 = 3.445838616e-07 wa0 = 1.277474911e-06 pa0 = -6.245191596e-13
+ ags = -4.184799672e+00 lags = 2.656910516e-06 wags = 3.041097154e-06 pags = -1.486701166e-12
+ a1 = 0.0
+ a2 = 6.945708973e+00 la2 = -2.930397677e-06 wa2 = -4.692809993e-06 pa2 = 2.294174021e-12
+ b0 = -3.145420887e-06 lb0 = 1.537701909e-12 wb0 = 2.502566057e-12 pb0 = -1.223429468e-18
+ b1 = -2.785872588e-07 lb1 = 1.361929532e-13 wb1 = 2.216501521e-13 pb1 = -1.083581098e-19
+ keta = -3.630914091e-01 lketa = 1.588449574e-07 wketa = 2.970258531e-07 pketa = -1.452070288e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.787427606e+00 lpclm = -3.289218088e-06 wpclm = -4.177874586e-06 ppclm = 2.042437549e-12
+ pdiblc1 = -1.012314940e+01 lpdiblc1 = 4.956513295e-06 wpdiblc1 = 8.103460008e-06 ppdiblc1 = -3.961538494e-12
+ pdiblc2 = 7.533057929e-04 lpdiblc2 = -3.197073994e-10
+ pdiblcb = 5.883813445e+00 lpdiblcb = -2.893755443e-06 wpdiblcb = -4.693044645e-06 ppdiblcb = 2.294288736e-12
+ drout = 8.812351559e+00 ldrout = -3.837722837e-06 wdrout = -6.186243096e-06 pdrout = 3.024268662e-12
+ pscbe1 = 4.190874397e+08 lpscbe1 = 1.611344822e+02 wpscbe1 = 3.214205268e+02 ppscbe1 = -1.571328529e-4
+ pscbe2 = 4.005175368e-09 lpscbe2 = 5.211869235e-15 wpscbe2 = -1.557011422e-16 ppscbe2 = 7.611761738e-23
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.193336930e+01 lbeta0 = -1.623331415e-05 wbeta0 = -2.808618036e-05 pbeta0 = 1.373049099e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.040850596e-08 lagidl = 9.977106307e-15 wagidl = 1.703690092e-14 pagidl = -8.328829752e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.254810687e-01 lkt1 = -5.298728500e-8
+ kt2 = -6.206186670e-02 lkt2 = 1.335240081e-8
+ at = 3.793635449e+05 lat = -1.666022485e-01 wat = -2.346522322e-01 pat = 1.147144368e-7
+ ute = -1.875821105e+00 lute = 8.184494349e-7
+ ua1 = -3.292299871e-09 lua1 = 2.830042980e-15 pua1 = -2.481541838e-36
+ ub1 = 5.214699782e-18 lub1 = -3.681876117e-24 wub1 = -9.386089290e-25 pub1 = 4.588577471e-31
+ uc1 = 3.136276955e-10 luc1 = -2.439630433e-16 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.141 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.809317576e-01 lvth0 = -1.208276190e-8
+ k1 = 4.446623754e-01 lk1 = 3.181784882e-8
+ k2 = 1.132757422e-02 lk2 = -5.805984424e-09 wk2 = 1.734723476e-24 pk2 = 4.336808690e-31
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.244403898e-01 ldsub = 2.171402925e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.700309796e-01 lvoff = -1.848941181e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.825934693e-01 lnfactor = 5.361094594e-7
+ eta0 = 4.169452362e-01 leta0 = 1.745059157e-8
+ etab = -1.210426333e-03 letab = 2.719825911e-10 petab = -4.336808690e-31
+ u0 = 4.591262030e-03 lu0 = 8.044064145e-10
+ ua = -1.330850367e-09 lua = 6.367127645e-17
+ ub = 7.875179014e-19 lub = 2.193322321e-25
+ uc = -6.000952568e-11 luc = 1.409804193e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.833766079e+04 lvsat = -2.582274881e-3
+ a0 = 8.732071908e-01 la0 = -6.153539006e-8
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 1.100021230e+00 la2 = -7.261631000e-8
+ b0 = 1.715100723e-16 lb0 = -4.096861098e-23
+ b1 = 7.130458861e-20 lb1 = -1.703252708e-26
+ keta = -4.438001254e-02 lketa = 3.036516966e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.930264200e-01 lpclm = 2.699774716e-07 wpclm = -2.220446049e-22 ppclm = 5.551115123e-29
+ pdiblc1 = -3.561786926e-01 lpdiblc1 = 1.817343246e-07 wpdiblc1 = -3.330669074e-22 ppdiblc1 = 2.081668171e-28
+ pdiblc2 = -8.000440691e-03 lpdiblc2 = 3.959736644e-09 wpdiblc2 = 2.602085214e-24 ppdiblc2 = 1.951563910e-30
+ pdiblcb = 2.058549522e-01 lpdiblcb = -1.179718745e-07 wpdiblcb = -2.220446049e-22 ppdiblcb = 2.775557562e-29
+ drout = 1.376341573e+00 ldrout = -2.024806355e-7
+ pscbe1 = 6.996965507e+08 lpscbe1 = 2.395310605e+1
+ pscbe2 = 2.022856548e-08 lpscbe2 = -2.719259489e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.553332902e+00 lbeta0 = 8.518424213e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.492459760e-12 lagidl = 7.296188029e-19
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.443546811e-01 lkt1 = 5.126457872e-9
+ kt2 = -1.748919269e-02 lkt2 = -8.437842332e-9
+ at = 1.056349506e+04 lat = 1.369303193e-2
+ ute = 4.030997005e-01 lute = -2.956465794e-7
+ ua1 = 4.600244176e-09 lua1 = -1.028385029e-15
+ ub1 = -4.368480081e-18 lub1 = 1.003053022e-24 wub1 = 6.162975822e-39
+ uc1 = -2.690313562e-10 luc1 = 4.088148730e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.142 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.126011471e+00 lvth0 = 2.257242935e-08 wvth0 = 2.156533171e-07 pvth0 = -5.151310785e-14
+ k1 = -1.995102558e+00 lk1 = 6.146044986e-07 wk1 = 1.030170672e-06 pk1 = -2.460768685e-13
+ k2 = 1.394589345e+00 lk2 = -3.362257236e-07 wk2 = -6.949977990e-07 pk2 = 1.660141242e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.029553202e+00 ldsub = -1.252864157e-06 wdsub = -3.280098685e-06 pdsub = 7.835171729e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.213650508e+00 lvoff = 2.307999848e-07 wvoff = 9.915767827e-07 pvoff = -2.368579461e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.186877128e+01 lnfactor = -2.064271835e-06 wnfactor = -7.724949905e-06 pnfactor = 1.845258784e-12
+ eta0 = 1.005205903e+01 leta0 = -2.284089039e-06 weta0 = -7.129681574e-06 peta0 = 1.703067038e-12
+ etab = 9.408004333e-01 letab = -2.247461515e-07 wetab = -7.001321498e-07 petab = 1.672405666e-13
+ u0 = 1.562974471e-03 lu0 = 1.527773464e-09 wu0 = 1.206161293e-08 pu0 = -2.881157480e-15
+ ua = -6.465954509e-09 lua = 1.290293603e-15 wua = 5.759885299e-15 pua = -1.375863801e-21
+ ub = 8.708471314e-18 lub = -1.672745910e-24 wub = -5.865942153e-24 pub = 1.401197602e-30
+ uc = -4.463702374e-10 luc = 1.063880251e-16 wuc = 3.542868288e-16 puc = -8.462849481e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.761679342e+04 lvsat = 2.272706560e-02 wvsat = 1.124520058e-01 pvsat = -2.686141062e-8
+ a0 = -9.070193890e+00 la0 = 2.313644826e-06 wa0 = 6.751502883e-06 pa0 = -1.612731494e-12
+ ags = 2.122259350e+00 lags = -1.472984343e-07 wags = 7.489404652e-15 pags = -1.788993842e-21
+ a1 = 0.0
+ a2 = 4.574808674e+00 la2 = -9.026387868e-07 wa2 = -2.732414667e-06 pa2 = 6.526918915e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.489558726e-01 lketa = 1.235645527e-07 wketa = 3.513232980e-07 pketa = -8.392059619e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.306276543e-01 lpclm = 1.570222884e-09 wpclm = 3.445359515e-08 ppclm = -8.229930273e-15
+ pdiblc1 = 7.158198815e+00 lpdiblc1 = -1.613225031e-06 wpdiblc1 = -4.946468176e-06 ppdiblc1 = 1.181562853e-12
+ pdiblc2 = -6.656347226e-02 lpdiblc2 = 1.794868799e-08 wpdiblc2 = 6.922782106e-08 ppdiblc2 = -1.653644962e-14
+ pdiblcb = -2.512532612e+01 lpdiblcb = 5.932887348e-06 wpdiblcb = 2.005006330e-05 ppdiblcb = -4.789358620e-12
+ drout = -6.083463697e-01 ldrout = 2.716017735e-07 wdrout = 3.383973521e-12 pdrout = -8.083297542e-19
+ pscbe1 = 7.999088715e+08 lpscbe1 = 1.538896829e-02 wpscbe1 = 1.012386322e-06 ppscbe1 = -2.418289185e-13
+ pscbe2 = -6.099503773e-08 lpscbe2 = 1.668262261e-14 wpscbe2 = 5.871176260e-14 ppscbe2 = -1.402447873e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033939091e+01 lbeta0 = -3.414514355e-07 wbeta0 = -6.571410038e-08 pbeta0 = 1.569712716e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.720009864e-08 lagidl = -8.885614448e-15 wagidl = -2.959555969e-14 pagidl = 7.069491343e-21
+ bgidl = 1.818113535e+09 lbgidl = -1.381548250e+02 wbgidl = 3.757583618e-06 pbgidl = -8.975744247e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.151191040e+00 lkt1 = 3.889514590e-07 wkt1 = 1.328849399e-06 pkt1 = -3.174222559e-13
+ kt2 = 1.552549457e+00 lkt2 = -3.834729746e-07 wkt2 = -1.200640066e-06 pkt2 = 2.867968925e-13
+ at = -6.261514054e+05 lat = 1.657851202e-01 wat = 6.067231435e-01 pat = -1.449279573e-7
+ ute = -1.702407539e+01 lute = 3.867182733e-06 wute = 1.143926410e-05 pute = -2.732497016e-12
+ ua1 = -1.377535434e-08 lua1 = 3.360994189e-15 wua1 = 1.039236170e-14 pua1 = -2.482423440e-21
+ ub1 = 1.239997046e-17 lub1 = -3.002426759e-24 wub1 = -9.471684215e-24 pub1 = 2.262501209e-30
+ uc1 = -5.240397428e-10 luc1 = 1.017953406e-16 wuc1 = 1.943816211e-16 puc1 = -4.643193783e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.143 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 6.483885964e-02 lvth0 = -1.964985743e-07 wvth0 = -8.658316030e-07 pvth0 = 1.443167133e-13
+ k1 = 3.720798198e+00 lk1 = -3.859382602e-07 wk1 = -2.029890744e-06 pk1 = 2.979243967e-13
+ k2 = -2.409003659e+00 lk2 = 3.369005489e-07 wk2 = 1.679760406e-06 pk2 = -2.586696819e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -8.000848692e+00 ldsub = 1.228841869e-06 wdsub = 6.463245402e-06 pdsub = -9.486021818e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 2.151630271e+00 lvoff = -3.714703144e-07 wvoff = -1.953126135e-06 pvoff = 2.866296961e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -1.592510396e+01 lnfactor = 2.893967257e-06 wnfactor = 1.521597346e-05 pnfactor = -2.233010003e-12
+ eta0 = -1.784372389e+01 leta0 = 2.670962820e-06 weta0 = 1.404345731e-05 peta0 = -2.060937969e-12
+ etab = -1.801253074e+00 letab = 2.622943291e-07 wetab = 1.379569570e-06 petab = -2.024776258e-13
+ u0 = 4.341176774e-02 lu0 = -6.096862079e-09 wu0 = -2.994303157e-08 pu0 = 4.636202107e-15
+ ua = 1.278400471e-08 lua = -2.157803552e-15 wua = -1.134535263e-14 pua = 1.664979728e-21
+ ub = -1.302000824e-17 lub = 2.197532670e-24 wub = 1.155424415e-23 pub = -1.695635049e-30
+ uc = 8.977215665e-10 luc = -1.327283260e-16 wuc = -6.981012433e-16 puc = 1.024593972e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.390200528e+05 lvsat = -4.127311056e-02 wvsat = -2.189225160e-01 pvsat = 3.202705626e-8
+ a0 = 1.823837799e+01 la0 = -2.529286762e-06 wa0 = -1.329854943e-05 pa0 = 1.951619415e-12
+ ags = 1.250000079e+00 lags = -1.228589142e-14 wags = -1.923450554e-14 pags = 2.998081783e-21
+ a1 = 0.0
+ a2 = -6.277752155e+00 la2 = 1.023658812e-06 wa2 = 5.384061670e-06 pa2 = -7.902116248e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 8.908599478e-01 lketa = -1.316148749e-07 wketa = -6.920079252e-07 pketa = 1.015551629e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.093695618e-01 lpclm = -1.290746246e-08 wpclm = -6.788850981e-08 ppclm = 9.963896660e-15
+ pdiblc1 = -1.236484697e+01 lpdiblc1 = 1.853121490e-06 wpdiblc1 = 9.746724286e-06 ppdiblc1 = -1.430513897e-12
+ pdiblc2 = 1.792574833e-01 lpdiblc2 = -2.593517378e-08 wpdiblc2 = -1.364093079e-07 ppdiblc2 = 2.002061315e-14
+ pdiblcb = 5.041997754e+01 lpdiblcb = -7.511459495e-06 wpdiblcb = -3.950746244e-05 ppdiblcb = 5.798458010e-12
+ drout = 1.000011818e+00 ldrout = -1.842213134e-12 wdrout = -8.690815633e-12 pdrout = 1.354637433e-18
+ pscbe1 = 8.000000039e+08 lpscbe1 = -6.168899536e-07 wpscbe1 = -2.600036621e-06 ppscbe1 = 4.052677155e-13
+ pscbe2 = 1.561327559e-07 lpscbe2 = -2.199549489e-14 wpscbe2 = -1.156880607e-13 ppscbe2 = 1.697938402e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.184954496e+00 lbeta0 = 2.462003450e-08 wbeta0 = 1.294897247e-07 pbeta0 = -1.900519131e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.555720624e-08 lagidl = 1.489547852e-14 wagidl = 7.601580889e-14 pagidl = -1.184881402e-20
+ bgidl = 1.000000282e+09 lbgidl = -4.388798332e-05 wbgidl = -9.650329590e-06 pbgidl = 1.504196167e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.830400378e+00 lkt1 = -4.978215236e-07 wkt1 = -2.617458700e-06 pkt1 = 3.841234006e-13
+ kt2 = -3.138249688e+00 lkt2 = 4.498019627e-07 wkt2 = 2.365789776e-06 pkt2 = -3.472238216e-13
+ at = 1.578477725e+06 lat = -2.272998486e-01 wat = -1.195512013e+00 pat = 1.754637164e-7
+ ute = 2.893299129e+01 lute = -4.285551235e-06 wute = -2.254039350e-05 pute = 3.308223781e-12
+ ua1 = 2.707408995e-08 lua1 = -3.893343580e-15 wua1 = -2.047752921e-14 pua1 = 3.005459716e-21
+ ub1 = -2.447045059e-17 lub1 = 3.548426641e-24 wub1 = 1.866339365e-23 pub1 = -2.739201632e-30
+ uc1 = 4.705542467e-10 luc1 = -7.282219343e-17 wuc1 = -3.830174561e-16 puc1 = 5.621496476e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.144 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.145 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108623478e+00 lvth0 = 3.532668562e-7
+ k1 = 4.171052081e-01 lk1 = 2.908460917e-7
+ k2 = 2.159455618e-02 lk2 = -4.690448662e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 2.541098842e-27 pcit = 2.710505431e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.807199248e-01 lvoff = 2.151443021e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.403205388e+00 lnfactor = -5.131826301e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.149534990e-02 lu0 = -1.176644632e-8
+ ua = -9.044296180e-10 lua = 2.075453526e-15
+ ub = 1.700362603e-18 lub = -5.753769297e-24
+ uc = -1.046578370e-10 luc = -2.009187197e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.286628951e+04 lvsat = -2.540643246e-1
+ a0 = 1.625827411e+00 la0 = -3.234747073e-6
+ ags = 1.127460711e-01 lags = 1.087252350e-8
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-06 wa2 = 1.776356839e-21
+ b0 = -2.227955321e-07 lb0 = 2.397975426e-12
+ b1 = 3.393294966e-09 lb1 = -2.149792907e-14
+ keta = 3.416681995e-02 lketa = -2.159909532e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 wpclm = -5.551115123e-23 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.906905271e-03 lpdiblc2 = -1.258792035e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.865952071e-09 lpscbe2 = 2.388016187e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.797495750e+01 lbeta0 = -3.592990887e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.808012713e-09 lagidl = -1.814500294e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443649873e-01 lkt1 = 1.222316870e-7
+ kt2 = -6.519461656e-02 lkt2 = 1.328983321e-7
+ at = 7.713361212e+04 lat = -1.228038641e-01 wat = -1.164153218e-16
+ ute = 5.595779957e-01 lute = -1.284400824e-05 pute = 3.552713679e-27
+ ua1 = 3.768264800e-09 lua1 = -3.354261913e-14 wua1 = -3.308722450e-30 pua1 = 2.646977960e-35
+ ub1 = -2.642787222e-18 lub1 = 2.826200788e-23
+ uc1 = -9.417115820e-11 luc1 = 1.286926591e-15 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.146 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.068784975e+00 lvth0 = 3.500223376e-8
+ k1 = 4.603509166e-01 lk1 = -5.463825109e-8
+ k2 = 1.538364979e-02 lk2 = 2.713637080e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.682810246e-01 lvoff = 1.157715452e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.131821908e+00 lnfactor = 5.025091038e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.814547492e-03 lu0 = 9.650135606e-9
+ ua = -8.481377777e-10 lua = 1.625745332e-15
+ ub = 1.054996270e-18 lub = -5.980215607e-25
+ uc = -1.070085284e-10 luc = -1.312504100e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342054363e+04 lvsat = -1.882608877e-2
+ a0 = 1.169648264e+00 la0 = 4.096088288e-7
+ ags = 4.536500838e-02 lags = 5.491710742e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 5.989974384e-08 lb0 = 1.395596165e-13
+ b1 = -9.045963073e-10 lb1 = 1.283736559e-14 pb1 = -6.617444900e-36
+ keta = 7.536869066e-03 lketa = -3.247737421e-09 wketa = -1.387778781e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.061808156e-01 lpclm = 4.371028699e-06 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.327209668e-04 lpdiblc2 = 7.869204170e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461096001e-08 lpscbe2 = -2.201595970e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.997217500e-10 lalpha0 = -7.966640969e-16
+ alpha1 = 1.997217500e-10 lalpha1 = -7.966640969e-16
+ beta0 = -2.392487250e+01 lbeta0 = 2.150993062e-04 pbeta0 = -2.842170943e-26
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.932747516e-10 lagidl = -1.250636281e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.139217330e-01 lkt1 = -1.209755144e-7
+ kt2 = -3.860015032e-02 lkt2 = -7.956140140e-8
+ at = 2.264263863e+04 lat = 3.125174394e-1
+ ute = -1.910932237e+00 lute = 6.892576840e-6
+ ua1 = -2.943994399e-09 lua1 = 2.008074701e-14 wua1 = -1.654361225e-30 pua1 = -6.617444900e-36
+ ub1 = 2.913039917e-18 lub1 = -1.612277288e-23
+ uc1 = 5.506278879e-10 luc1 = -3.864289165e-15 puc1 = -2.481541838e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.147 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.063486545e+00 lvth0 = 1.386748510e-8
+ k1 = 3.863911154e-01 lk1 = 2.403777808e-7
+ k2 = 3.756574616e-02 lk2 = -8.576786165e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.583304901e-01 ldsub = -1.190001542e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.481840352e-01 lvoff = 3.560726699e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.206074825e+00 lnfactor = 7.400358035e-7
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391132325e-01 letab = 2.756836997e-7
+ u0 = 1.129796699e-02 lu0 = -2.559019068e-10
+ ua = -3.948101738e-10 lua = -1.825195469e-16
+ ub = 9.047694627e-19 lub = 1.213642946e-27
+ uc = -1.333555795e-10 luc = 1.037824576e-16 wuc = 2.067951531e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.345823238e+04 lvsat = -9.875382428e-2
+ a0 = 1.398566000e+00 la0 = -5.035142625e-7
+ ags = -4.042771799e-02 lags = 8.913871067e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 7.545275680e-08 lb0 = 7.752066969e-14
+ b1 = 6.234956092e-09 lb1 = -1.564138079e-14
+ keta = 2.253544784e-02 lketa = -6.307511832e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.074223900e-01 lpclm = 3.278972801e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.187393462e-04 lpdiblc2 = 4.491728403e-11
+ pdiblcb = -4.238870000e-01 lpdiblcb = 7.933343877e-07 ppdiblcb = 8.881784197e-28
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.718970657e-09 lpscbe2 = 1.486419869e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.944350000e-11 lalpha0 = 3.966671938e-16
+ alpha1 = -9.944350000e-11 lalpha1 = 3.966671938e-16
+ beta0 = 5.429614004e+01 lbeta0 = -9.691414411e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.573122120e-11 lagidl = 1.776939874e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356779703e-01 lkt1 = -3.419271211e-8
+ kt2 = -6.313133978e-02 lkt2 = 1.829032431e-8
+ at = 1.615988244e+05 lat = -2.417607213e-1
+ ute = -9.311290905e-02 lute = -3.584681431e-7
+ ua1 = 2.873317563e-09 lua1 = -3.123754152e-15
+ ub1 = -1.891532201e-18 lub1 = 3.042040710e-24 wub1 = -3.081487911e-39
+ uc1 = -8.692813487e-10 luc1 = 1.799544192e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.148 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.081021165e+00 lvth0 = 4.874156567e-8
+ k1 = 5.064919019e-01 lk1 = 1.512929702e-9
+ k2 = -5.250837621e-03 lk2 = -6.112426770e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000199e-01 ldsub = -1.966733887e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.231624387e-01 lvoff = -1.415743548e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.405520147e+00 lnfactor = 3.433649873e-7
+ eta0 = -4.835518650e-01 leta0 = 9.627162327e-07 weta0 = 4.180683577e-22 peta0 = -7.372574773e-28
+ etab = 2.386594872e-04 letab = -1.469097694e-9
+ u0 = 1.277578903e-02 lu0 = -3.195097838e-9
+ ua = -2.787126111e-10 lua = -4.134225064e-16
+ ub = 8.338866336e-19 lub = 1.421903751e-25
+ uc = -1.183445084e-10 luc = 7.392738859e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.599790864e+04 lvsat = 3.541598979e-2
+ a0 = 1.034813481e+00 la0 = 2.199422095e-7
+ ags = 2.529917783e-01 lags = 3.078138731e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.221234086e-07 lb0 = -1.530118956e-14
+ b1 = -1.258163080e-08 lb1 = 2.178236438e-14 pb1 = 3.308722450e-36
+ keta = -1.722971284e-02 lketa = 1.601261680e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.149196182e-01 lpclm = -2.836747322e-7
+ pdiblc1 = 3.955978546e-01 lpdiblc1 = -1.113340513e-8
+ pdiblc2 = 4.525213076e-04 lpdiblc2 = -2.227064540e-11
+ pdiblcb = 1.727740000e-01 lpdiblcb = -3.933467754e-7
+ drout = 3.855974777e-01 ldrout = 3.468639446e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.759262277e-09 lpscbe2 = -5.825849256e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.674544110e+00 lbeta0 = 1.776759381e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.258387184e-10 lagidl = 7.992711679e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.269668075e-01 lkt1 = -5.151808255e-8
+ kt2 = -5.925098613e-02 lkt2 = 1.057280534e-8
+ at = 2.845269774e+04 lat = 2.304961559e-2
+ ute = 4.928361669e-01 lute = -1.523844682e-06 pute = 8.881784197e-28
+ ua1 = 3.016514543e-09 lua1 = -3.408554329e-15
+ ub1 = -1.565341614e-18 lub1 = 2.393290035e-24 pub1 = 7.703719778e-46
+ uc1 = 4.482619664e-12 luc1 = 6.174124785e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.149 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.131471245e+00 lvth0 = 9.863013585e-08 wvth0 = 5.535297701e-08 pvth0 = -5.473689837e-14
+ k1 = -3.293797507e-01 lk1 = 8.280813307e-07 wk1 = 6.231275013e-07 pk1 = -6.161920922e-13
+ k2 = 2.736935042e-01 lk2 = -2.764509339e-07 wk2 = -2.123264782e-07 pk2 = 2.099632845e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.802062121e+00 ldsub = -7.458118970e-06 wdsub = -5.667070156e-06 pdsub = 5.603995665e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -6.735997778e-01 lvoff = 4.312665359e-07 wvoff = 3.035818903e-07 pvoff = -3.002030238e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.789854678e+01 lnfactor = -3.475462426e-05 wnfactor = -2.571446220e-05 pnfactor = 2.542826023e-11
+ eta0 = -4.439393457e+00 leta0 = 4.874529308e-06 weta0 = 3.702699827e-06 peta0 = -3.661488778e-12
+ etab = -5.691544758e-03 letab = 4.395103378e-09 wetab = 2.881734220e-09 petab = -2.849660518e-15
+ u0 = 2.032741929e-01 lu0 = -1.915732545e-07 wu0 = -1.420373173e-07 pu0 = 1.404564420e-13
+ ua = 2.666685468e-08 lua = -2.705908563e-14 wua = -2.003563686e-14 pua = 1.981264022e-20
+ ub = 7.139574768e-18 lub = -6.093315450e-24 wub = -4.782893190e-24 pub = 4.729659589e-30
+ uc = -2.474564145e-10 luc = 2.016022792e-16 wuc = 1.429612030e-16 puc = -1.413700448e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.426952333e+05 lvsat = 2.912298771e-01 wvsat = 1.968145338e-01 pvsat = -1.946239880e-7
+ a0 = 5.855761333e+00 la0 = -4.547348493e-06 wa0 = -3.057038060e-06 pa0 = 3.023013226e-12
+ ags = -1.061952935e-01 lags = 6.630031928e-07 wags = -4.920881480e-16 pags = 4.866116399e-22
+ a1 = 0.0
+ a2 = -4.480007950e+00 la2 = 5.221241461e-06 wa2 = 3.826455911e-06 pa2 = -3.783867457e-12
+ b0 = 2.109259699e-07 lb0 = -1.031153784e-13 wb0 = 7.306542202e-22 pb0 = -7.225219627e-28
+ b1 = 1.868153427e-08 lb1 = -9.132841656e-15 wb1 = 3.037671907e-25 pb1 = -3.003790589e-31
+ keta = -2.464260546e-02 lketa = 2.334300392e-08 wketa = 4.467097925e-08 pketa = -4.417379126e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.354807759e+00 lpclm = -4.674146918e-06 wpclm = -3.109681710e-06 ppclm = 3.075070953e-12
+ pdiblc1 = 1.351662203e+00 lpdiblc1 = -9.565567569e-07 wpdiblc1 = -4.524119689e-07 ppdiblc1 = 4.473766237e-13
+ pdiblc2 = 8.622179337e-03 lpdiblc2 = -8.101000381e-09 wpdiblc2 = -5.867205230e-09 ppdiblc2 = 5.801903235e-15
+ pdiblcb = -2.527982441e+00 lpdiblcb = 2.277350246e-06 wpdiblcb = 1.578975427e-06 ppdiblcb = -1.561401431e-12
+ drout = -4.514177379e+00 ldrout = 5.192104307e-06 wdrout = 3.750310063e-06 pdrout = -3.708569112e-12
+ pscbe1 = -5.969729043e+09 lpscbe1 = 6.694381959e+03 wpscbe1 = 5.085062650e+03 ppscbe1 = -5.028465903e-3
+ pscbe2 = 7.133571335e-07 lpscbe2 = -6.963494119e-13 wpscbe2 = -5.290641269e-13 ppscbe2 = 5.231756431e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.075903012e+00 lbeta0 = 5.335347604e-06 wbeta0 = 2.378045367e-06 pbeta0 = -2.351577723e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.264582053e-08 lagidl = -1.128470224e-14 wagidl = -7.609132103e-15 pagidl = 7.524442463e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.330220297e-01 lkt1 = -6.052742439e-07 wkt1 = -4.164321972e-07 pkt1 = 4.117973069e-13
+ kt2 = -3.390872373e-01 lkt2 = 2.872944791e-07 wkt2 = 2.065562109e-07 pkt2 = -2.042572403e-13
+ at = 5.275063766e+05 lat = -4.704495958e-01 wat = -3.451107867e-01 pat = 3.412697036e-7
+ ute = -2.288591904e+00 lute = 1.226626094e-06 wute = 3.077709884e-07 pute = -3.043454973e-13
+ ua1 = -1.257732369e-08 lua1 = 1.201172448e-14 wua1 = 6.923118031e-15 pua1 = -6.846063727e-21
+ ub1 = 2.015916203e-17 lub1 = -1.908941988e-23 wub1 = -1.208152876e-23 pub1 = 1.194706134e-29
+ uc1 = 1.632649380e-09 luc1 = -1.548304017e-15 wuc1 = -9.834915867e-16 puc1 = 9.725453254e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.150 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.324571230e-01 lvth0 = -4.754889788e-08 wvth0 = -1.107059540e-07 pvth0 = 2.644433124e-14
+ k1 = 2.116092406e+00 lk1 = -3.674366427e-07 wk1 = -1.246255003e-06 pk1 = 2.976929325e-13
+ k2 = -5.582008952e-01 lk2 = 1.302372811e-07 wk2 = 4.246529564e-07 pk2 = -1.014368517e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.532536031e+01 ldsub = 3.848184034e-06 wdsub = 1.133414031e-05 pdsub = -2.707386096e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 6.442740980e-01 lvoff = -2.130024657e-07 wvoff = -6.071637805e-07 pvoff = 1.450332123e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -6.799193302e+01 lnfactor = 1.701205460e-05 wnfactor = 5.142892439e-05 pnfactor = -1.228482717e-11
+ eta0 = 1.034878691e+01 leta0 = -2.354968430e-06 weta0 = -7.405399655e-06 peta0 = 1.768927816e-12
+ etab = 6.519319356e-03 letab = -1.574421762e-09 wetab = -5.763468440e-09 petab = 1.376719706e-15
+ u0 = -3.763988839e-01 lu0 = 9.181152258e-08 wu0 = 2.840746346e-07 pu0 = -6.785690797e-14
+ ua = -5.507292573e-08 lua = 1.290104082e-14 wua = 4.007127372e-14 pua = -9.571825153e-21
+ ub = -1.204175267e-17 lub = 3.283860093e-24 wub = 9.565786380e-24 pub = -2.284979393e-30
+ uc = 3.234587812e-10 luc = -7.750103253e-17 wuc = -2.859224059e-16 puc = 6.829828510e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.162580649e+05 lvsat = -1.286866218e-01 wvsat = -3.936290675e-01 pvsat = 9.402617536e-8
+ a0 = -7.326760246e+00 la0 = 1.897190832e-06 wa0 = 6.114076120e-06 pa0 = -1.460469363e-12
+ ags = 1.005767372e+00 lags = 1.193980046e-07 wags = 9.841762960e-16 pags = -2.350910577e-22
+ a1 = 0.0
+ a2 = 1.136381686e+01 la2 = -2.524329171e-06 wa2 = -7.652911822e-06 pa2 = 1.828051047e-12
+ b0 = 2.131361386e-15 lb0 = -5.091182942e-22 wb0 = -1.461308256e-21 pb0 = 3.490627031e-28
+ b1 = 8.861044995e-19 lb1 = -2.116637818e-25 wb1 = -6.075327392e-25 pb1 = 1.451213454e-31
+ keta = 7.544204007e-02 lketa = -2.558537674e-08 wketa = -8.934195851e-08 pketa = 2.134111363e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -8.834201198e+00 lpclm = 2.262433891e-06 wpclm = 6.219363421e-06 ppclm = -1.485619340e-12
+ pdiblc1 = -1.569694305e+00 lpdiblc1 = 4.716067989e-07 wpdiblc1 = 9.048239377e-07 ppdiblc1 = -2.161352940e-13
+ pdiblc2 = -2.373818778e-02 lpdiblc2 = 7.719012291e-09 wpdiblc2 = 1.173441046e-08 ppdiblc2 = -2.802998626e-15
+ pdiblcb = 4.441179090e+00 lpdiblcb = -1.129663751e-06 wpdiblcb = -3.157950854e-06 ppdiblcb = 7.543397206e-13
+ drout = 1.143588934e+01 ldrout = -2.605404811e-06 wdrout = -7.500620127e-06 pdrout = 1.791673130e-12
+ pscbe1 = 1.433948360e+10 lpscbe1 = -3.234182827e+03 wpscbe1 = -1.017012530e+04 ppscbe1 = 2.429337831e-3
+ pscbe2 = -1.398892992e-06 lpscbe2 = 3.362663069e-13 wpscbe2 = 1.058128254e-12 ppscbe2 = -2.527550960e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.493202175e+01 lbeta0 = -1.438493163e-06 wbeta0 = -4.756090735e-06 pbeta0 = 1.136087394e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.041165231e-08 lagidl = 4.876104502e-15 wagidl = 1.521826421e-14 pagidl = -3.635186771e-21
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.661360878e+00 lkt1 = 2.719457281e-07 wkt1 = 8.328643945e-07 pkt1 = -1.989463179e-13
+ kt2 = 5.365615486e-01 lkt2 = -1.407839429e-07 wkt2 = -4.131124218e-07 pkt2 = 9.868016420e-14
+ at = -9.151355499e+05 lat = 2.348147628e-01 wat = 6.902215733e-01 pat = -1.648732272e-7
+ ute = 1.228641298e+00 lute = -4.928437007e-07 wute = -6.155419767e-07 pute = 1.470345120e-13
+ ua1 = 2.317029182e-08 lua1 = -5.464212308e-15 wua1 = -1.384623606e-14 pua1 = 3.307450408e-21
+ ub1 = -3.677505811e-17 lub1 = 8.744012315e-24 wub1 = 2.416305752e-23 pub1 = -5.771829550e-30
+ uc1 = -2.907074726e-09 luc1 = 6.710309070e-16 wuc1 = 1.966983173e-15 puc1 = -4.698532706e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.151 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.367854064e-01 lvth0 = -4.651500081e-8
+ k1 = -6.134766510e-01 lk1 = 2.845755181e-7
+ k2 = 4.624846070e-01 lk2 = -1.135738648e-07 wk2 = -1.110223025e-22 pk2 = 2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.630409017e+00 ldsub = -2.020405853e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.162147361e-01 lvoff = -8.686492591e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.508360907e+00 lnfactor = 4.105193916e-7
+ eta0 = 4.900000007e-01 leta0 = -5.141975734e-17
+ etab = 1.809698392e-03 letab = -4.494346021e-10 wetab = 4.336808690e-25 petab = -1.626303259e-31
+ u0 = 1.773955312e-02 lu0 = -2.336325879e-9
+ ua = 1.258985607e-09 lua = -5.549628425e-16
+ ub = 8.412917613e-19 lub = 2.064872702e-25
+ uc = 2.878584554e-11 luc = -7.112508390e-18 wuc = 6.462348536e-33 puc = 3.231174268e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.331995797e+05 lvsat = -1.329844146e-2
+ a0 = -1.533380897e-02 la0 = 1.507103985e-7
+ ags = 2.122259360e+00 lags = -1.472984367e-7
+ a1 = 0.0
+ a2 = 9.101975611e-01 la2 = -2.727313031e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.777436513e-02 lketa = 1.101342597e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.768355118e-01 lpclm = -9.467448044e-9
+ pdiblc1 = 5.241829513e-01 lpdiblc1 = -2.855766128e-8
+ pdiblc2 = 2.628226065e-02 lpdiblc2 = -4.229372224e-09 wpdiblc2 = 2.775557562e-23
+ pdiblcb = 1.765059758e+00 lpdiblcb = -4.904191263e-07 ppdiblcb = -4.440892099e-28
+ drout = -6.083418313e-01 ldrout = 2.716006894e-7
+ pscbe1 = 7.999088729e+08 lpscbe1 = 1.538864396e-2
+ pscbe2 = 1.774695567e-08 lpscbe2 = -2.126477355e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025125765e+01 lbeta0 = -3.203990428e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.492345636e-09 lagidl = 5.957197170e-16 wagidl = 1.421716678e-30 pagidl = 2.391068958e-37
+ bgidl = 1.818113540e+09 lbgidl = -1.381548262e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.689885319e-01 lkt1 = -3.676325419e-8
+ kt2 = -5.770354749e-02 lkt2 = 1.168160598e-9
+ at = 1.875627065e+05 lat = -2.858676971e-2
+ ute = -1.682167421e+00 lute = 2.024611778e-7
+ ua1 = 1.624877580e-10 lua1 = 3.166184703e-17
+ ub1 = -3.030938486e-19 lub1 = 3.195421259e-26
+ uc1 = -2.633424711e-10 luc1 = 3.952258331e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.152 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.152383921e-01 lvth0 = -3.661557013e-08 wvth0 = -1.350644425e-07 pvth0 = 2.510442792e-14
+ k1 = 1.606404155e-01 lk1 = 1.693383555e-07 wk1 = 6.246412223e-07 pk1 = -1.161020640e-13
+ k2 = 4.596853226e-01 lk2 = -1.244869467e-07 wk2 = -4.591972097e-07 pk2 = 8.535098538e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.334815479e+00 ldsub = -5.391778692e-07 wdsub = -1.988875188e-06 pdsub = 3.696722312e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.263767247e+00 lvoff = 1.608877068e-07 wvoff = 5.934693943e-07 pvoff = -1.103081563e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.068279278e+01 lnfactor = -1.253405621e-06 wnfactor = -4.623459717e-06 pnfactor = 8.593624576e-13
+ eta0 = 6.713823862e+00 leta0 = -1.156822141e-06 weta0 = -4.267190562e-06 peta0 = 7.931427097e-13
+ etab = 6.183274690e-01 letab = -1.150868368e-07 wetab = -4.245229134e-07 petab = 7.890607392e-14
+ u0 = -4.187701093e-03 lu0 = 1.504096913e-09 wu0 = 5.548179579e-09 pu0 = -1.031240138e-15
+ ua = -7.055403364e-09 lua = 9.345649958e-16 wua = 3.447346496e-15 pua = -6.407582933e-22
+ ub = 7.184684656e-18 lub = -9.517722683e-25 wub = -3.510819380e-24 pub = 6.525559982e-31
+ uc = -3.266551770e-10 luc = 5.823730427e-17 wuc = 2.148209930e-16 puc = -3.992877797e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.789709698e+04 lvsat = 2.088195499e-02 wvsat = 7.702764312e-02 pvsat = -1.431712803e-8
+ a0 = -5.016567780e+00 la0 = 1.095461645e-06 wa0 = 4.040849743e-06 pa0 = -7.510727417e-13
+ ags = 1.250000052e+00 lags = -8.145683239e-15 wags = 4.785505325e-16 pags = -8.894573966e-23
+ a1 = 0.0
+ a2 = 3.165175715e+00 la2 = -4.491514827e-07 wa2 = -1.656793094e-06 pa2 = 3.079481325e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.192415940e-01 lketa = 5.700365207e-08 wketa = 2.102704067e-07 pketa = -3.908296049e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.903016768e-01 lpclm = 5.663515886e-09 wpclm = 2.089112475e-08 ppclm = -3.883033357e-15
+ pdiblc1 = 4.729608978e+00 lpdiblc1 = -8.130950725e-07 wpdiblc1 = -2.999278144e-06 ppdiblc1 = 5.574758287e-13
+ pdiblc2 = -5.998633668e-02 lpdiblc2 = 1.137960464e-08 wpdiblc2 = 4.197614767e-08 ppdiblc2 = -7.802106568e-15
+ pdiblcb = -1.887086035e+01 lpdiblcb = 3.295809265e-06 wpdiblcb = 1.215731069e-05 ppdiblcb = -2.259679337e-12
+ drout = 1.000000188e+00 ldrout = -3.018088357e-14 wdrout = -1.907957881e-14 pdrout = 3.546320571e-21
+ pscbe1 = 8.000000016e+08 lpscbe1 = -2.826652527e-07 wpscbe1 = -8.396453857e-07 ppscbe1 = 1.560640335e-13
+ pscbe2 = -4.676870923e-08 lpscbe2 = 9.650978605e-15 wpscbe2 = 3.559973552e-14 ppscbe2 = -6.616922840e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.412055214e+00 lbeta0 = -1.080078633e-08 wbeta0 = -3.984156649e-08 pbeta0 = 7.405351963e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.760675147e-08 lagidl = -1.237362886e-14 wagidl = -4.564282758e-14 pagidl = 8.483632363e-21
+ bgidl = 1.000000253e+09 lbgidl = -3.883447075e-05 wbgidl = 1.217955780e-05 pbgidl = -2.263813972e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.746702596e+00 lkt1 = 2.156115332e-07 wkt1 = 7.953299733e-07 pkt1 = -1.478279821e-13
+ kt2 = 1.011031791e+00 lkt2 = -1.973600790e-07 wkt2 = -7.280057794e-07 pkt2 = 1.353144342e-13
+ at = -5.182914647e+05 lat = 9.973253917e-02 wat = 3.678852243e-01 pat = -6.837882665e-8
+ ute = -1.059986113e+01 lute = 1.880374504e-06 wute = 6.936170982e-06 pute = -1.289226100e-12
+ ua1 = -8.840781778e-09 lua1 = 1.708286927e-15 wua1 = 6.301389280e-15 pua1 = -1.171239225e-21
+ ub1 = 8.262659774e-18 lub1 = -1.556945610e-24 wub1 = -5.743133568e-24 pub1 = 1.067476236e-30
+ uc1 = -2.012074926e-10 luc1 = 3.195225987e-17 wuc1 = 1.178628755e-16 puc1 = -2.190717267e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.153 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.154 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108623478e+00 lvth0 = 3.532668562e-7
+ k1 = 4.171052081e-01 lk1 = 2.908460917e-7
+ k2 = 2.159455618e-02 lk2 = -4.690448662e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = -2.032879073e-26 pcit = -1.084202172e-31
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.807199248e-01 lvoff = 2.151443021e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.403205388e+00 lnfactor = -5.131826301e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.149534990e-02 lu0 = -1.176644632e-8
+ ua = -9.044296180e-10 lua = 2.075453526e-15
+ ub = 1.700362603e-18 lub = -5.753769297e-24
+ uc = -1.046578370e-10 luc = -2.009187197e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.286628951e+04 lvsat = -2.540643246e-1
+ a0 = 1.625827411e+00 la0 = -3.234747073e-6
+ ags = 1.127460711e-01 lags = 1.087252350e-8
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = -2.227955321e-07 lb0 = 2.397975426e-12 pb0 = -1.355252716e-32
+ b1 = 3.393294966e-09 lb1 = -2.149792907e-14
+ keta = 3.416681995e-02 lketa = -2.159909532e-07 pketa = -1.776356839e-27
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.906905271e-03 lpdiblc2 = -1.258792035e-08 wpdiblc2 = -1.387778781e-23
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.865952071e-09 lpscbe2 = 2.388016187e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.797495750e+01 lbeta0 = -3.592990887e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.808012713e-09 lagidl = -1.814500294e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443649873e-01 lkt1 = 1.222316870e-7
+ kt2 = -6.519461656e-02 lkt2 = 1.328983321e-7
+ at = 7.713361212e+04 lat = -1.228038641e-1
+ ute = 5.595779957e-01 lute = -1.284400824e-05 wute = 8.881784197e-22 pute = -5.684341886e-26
+ ua1 = 3.768264800e-09 lua1 = -3.354261913e-14 pua1 = -2.117582368e-34
+ ub1 = -2.642787222e-18 lub1 = 2.826200788e-23 pub1 = 9.860761315e-44
+ uc1 = -9.417115820e-11 luc1 = 1.286926591e-15 puc1 = -6.617444900e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.155 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.068784975e+00 lvth0 = 3.500223376e-8
+ k1 = 4.603509166e-01 lk1 = -5.463825109e-8
+ k2 = 1.538364979e-02 lk2 = 2.713637080e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.682810246e-01 lvoff = 1.157715452e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.131821908e+00 lnfactor = 5.025091038e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.814547492e-03 lu0 = 9.650135606e-9
+ ua = -8.481377777e-10 lua = 1.625745332e-15
+ ub = 1.054996270e-18 lub = -5.980215607e-25
+ uc = -1.070085284e-10 luc = -1.312504100e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342054363e+04 lvsat = -1.882608877e-2
+ a0 = 1.169648264e+00 la0 = 4.096088288e-7
+ ags = 4.536500838e-02 lags = 5.491710742e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 5.989974383e-08 lb0 = 1.395596165e-13
+ b1 = -9.045963073e-10 lb1 = 1.283736559e-14
+ keta = 7.536869066e-03 lketa = -3.247737421e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.061808156e-01 lpclm = 4.371028699e-06 ppclm = -7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.327209668e-04 lpdiblc2 = 7.869204170e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461096001e-08 lpscbe2 = -2.201595970e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.997217500e-10 lalpha0 = -7.966640969e-16
+ alpha1 = 1.997217500e-10 lalpha1 = -7.966640969e-16
+ beta0 = -2.392487250e+01 lbeta0 = 2.150993062e-04 wbeta0 = -5.684341886e-20 pbeta0 = -6.821210263e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.932747516e-10 lagidl = -1.250636281e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.139217330e-01 lkt1 = -1.209755144e-7
+ kt2 = -3.860015032e-02 lkt2 = -7.956140140e-8
+ at = 2.264263863e+04 lat = 3.125174394e-1
+ ute = -1.910932237e+00 lute = 6.892576840e-6
+ ua1 = -2.943994399e-09 lua1 = 2.008074701e-14 wua1 = -1.323488980e-29 pua1 = 5.293955920e-35
+ ub1 = 2.913039917e-18 lub1 = -1.612277288e-23 wub1 = 1.232595164e-38 pub1 = -4.930380658e-44
+ uc1 = 5.506278879e-10 luc1 = -3.864289165e-15 wuc1 = -8.271806126e-31 puc1 = -6.617444900e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.156 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.063486545e+00 lvth0 = 1.386748510e-8
+ k1 = 3.863911154e-01 lk1 = 2.403777808e-7
+ k2 = 3.756574616e-02 lk2 = -8.576786165e-08 pk2 = -4.440892099e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.583304901e-01 ldsub = -1.190001542e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.481840352e-01 lvoff = 3.560726699e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.206074825e+00 lnfactor = 7.400358035e-7
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391132325e-01 letab = 2.756836997e-7
+ u0 = 1.129796699e-02 lu0 = -2.559019068e-10
+ ua = -3.948101738e-10 lua = -1.825195469e-16
+ ub = 9.047694627e-19 lub = 1.213642946e-27
+ uc = -1.333555795e-10 luc = 1.037824576e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.345823238e+04 lvsat = -9.875382428e-2
+ a0 = 1.398566000e+00 la0 = -5.035142625e-7
+ ags = -4.042771799e-02 lags = 8.913871067e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 7.545275680e-08 lb0 = 7.752066969e-14
+ b1 = 6.234956092e-09 lb1 = -1.564138079e-14 wb1 = -2.646977960e-29 pb1 = 5.293955920e-35
+ keta = 2.253544784e-02 lketa = -6.307511832e-08 wketa = 1.110223025e-22 pketa = 2.220446049e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.074223900e-01 lpclm = 3.278972801e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.187393462e-04 lpdiblc2 = 4.491728403e-11
+ pdiblcb = -4.238870000e-01 lpdiblcb = 7.933343877e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.718970657e-09 lpscbe2 = 1.486419869e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.944350000e-11 lalpha0 = 3.966671938e-16
+ alpha1 = -9.944350000e-11 lalpha1 = 3.966671938e-16
+ beta0 = 5.429614004e+01 lbeta0 = -9.691414411e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.573122120e-11 lagidl = 1.776939874e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356779703e-01 lkt1 = -3.419271211e-8
+ kt2 = -6.313133979e-02 lkt2 = 1.829032431e-8
+ at = 1.615988244e+05 lat = -2.417607213e-1
+ ute = -9.311290905e-02 lute = -3.584681431e-7
+ ua1 = 2.873317563e-09 lua1 = -3.123754152e-15
+ ub1 = -1.891532202e-18 lub1 = 3.042040710e-24
+ uc1 = -8.692813487e-10 luc1 = 1.799544192e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.157 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.081021165e+00 lvth0 = 4.874156567e-8
+ k1 = 5.064919019e-01 lk1 = 1.512929702e-9
+ k2 = -5.250837621e-03 lk2 = -6.112426770e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000199e-01 ldsub = -1.966733976e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.231624387e-01 lvoff = -1.415743548e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.405520147e+00 lnfactor = 3.433649873e-7
+ eta0 = -4.835518650e-01 leta0 = 9.627162327e-07 weta0 = 6.383782392e-22 peta0 = -1.991462550e-27
+ etab = 2.386594872e-04 letab = -1.469097694e-09 petab = 6.938893904e-30
+ u0 = 1.277578903e-02 lu0 = -3.195097838e-9
+ ua = -2.787126111e-10 lua = -4.134225064e-16
+ ub = 8.338866336e-19 lub = 1.421903751e-25
+ uc = -1.183445084e-10 luc = 7.392738859e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.599790864e+04 lvsat = 3.541598979e-2
+ a0 = 1.034813481e+00 la0 = 2.199422095e-7
+ ags = 2.529917783e-01 lags = 3.078138731e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.221234086e-07 lb0 = -1.530118956e-14
+ b1 = -1.258163080e-08 lb1 = 2.178236438e-14 wb1 = 2.646977960e-29 pb1 = -2.646977960e-35
+ keta = -1.722971284e-02 lketa = 1.601261680e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.149196182e-01 lpclm = -2.836747322e-7
+ pdiblc1 = 3.955978546e-01 lpdiblc1 = -1.113340513e-8
+ pdiblc2 = 4.525213076e-04 lpdiblc2 = -2.227064540e-11
+ pdiblcb = 1.727740000e-01 lpdiblcb = -3.933467754e-7
+ drout = 3.855974777e-01 ldrout = 3.468639446e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.759262277e-09 lpscbe2 = -5.825849256e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.674544110e+00 lbeta0 = 1.776759381e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.258387184e-10 lagidl = 7.992711679e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.269668075e-01 lkt1 = -5.151808255e-8
+ kt2 = -5.925098613e-02 lkt2 = 1.057280534e-8
+ at = 2.845269774e+04 lat = 2.304961559e-2
+ ute = 4.928361669e-01 lute = -1.523844682e-06 pute = -3.552713679e-27
+ ua1 = 3.016514543e-09 lua1 = -3.408554329e-15
+ ub1 = -1.565341614e-18 lub1 = 2.393290035e-24
+ uc1 = 4.482619664e-12 luc1 = 6.174124785e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.158 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.050737288e+00 lvth0 = 1.879474788e-8
+ k1 = 5.794701714e-01 lk1 = -7.065309168e-8
+ k2 = -3.599095491e-02 lk2 = 2.978673710e-08 wk2 = -1.110223025e-22 pk2 = -5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.635276000e-01 ldsub = 7.154747378e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.308165965e-01 lvoff = -6.588468460e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.932418197e-01 lnfactor = 2.333246657e-6
+ eta0 = 9.611039418e-01 leta0 = -4.658605549e-7
+ etab = -1.488450021e-03 letab = 2.387890846e-10
+ u0 = -3.891442511e-03 lu0 = 1.328662742e-8
+ ua = -2.555715282e-09 lua = 1.838237125e-15
+ ub = 1.635833473e-19 lub = 8.050331859e-25
+ uc = -3.894326448e-11 luc = -4.590119479e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.436459522e+04 lvsat = 7.365024437e-3
+ a0 = 1.396980751e+00 la0 = -1.381941390e-7
+ ags = -1.061952942e-01 lags = 6.630031935e-7
+ a1 = 0.0
+ a2 = 1.100991363e+00 la2 = -2.976413294e-7
+ b0 = 2.109259710e-07 lb0 = -1.031153794e-13
+ b1 = 1.868153427e-08 lb1 = -9.132841657e-15
+ keta = 4.051134126e-02 lketa = -4.108577937e-08 wketa = 8.326672685e-23 pketa = 1.387778781e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.192448538e-01 lpclm = -1.890648279e-7
+ pdiblc1 = 6.918059423e-01 lpdiblc1 = -3.040446968e-07 wpdiblc1 = 7.105427358e-21
+ pdiblc2 = 6.468668115e-05 lpdiblc2 = 3.612473816e-10
+ pdiblcb = -0.225
+ drout = 9.557609593e-01 ldrout = -2.169536175e-7
+ pscbe1 = 1.446985488e+09 lpscbe1 = -6.397845396e+2
+ pscbe2 = -5.829857018e-08 lpscbe2 = 6.671776386e-14 ppscbe2 = -1.588186776e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.544352635e+00 lbeta0 = 1.905501825e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.547675918e-09 lagidl = -3.100799834e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.743566677e-01 lkt1 = -4.655671468e-9
+ kt2 = -3.781888407e-02 lkt2 = -1.062075742e-8
+ at = 2.415206960e+04 lat = 2.730237773e-2
+ ute = -1.839698799e+00 lute = 7.827291698e-7
+ ua1 = -2.479750931e-09 lua1 = 2.026537710e-15 pua1 = 6.617444900e-36
+ ub1 = 2.537894393e-18 lub1 = -1.664276955e-24 pub1 = -6.162975822e-45
+ uc1 = 1.981977632e-10 luc1 = -1.298178461e-16 wuc1 = -8.271806126e-31 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.159 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.939250368e-01 lvth0 = -8.979057300e-9
+ k1 = 2.983925622e-01 lk1 = 6.675731910e-8
+ k2 = 6.116802299e-02 lk2 = -1.771137242e-08 pk2 = -1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.205819134e+00 ldsub = -1.006188000e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.412922644e-01 lvoff = -1.467228692e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.018676894e+00 lnfactor = -9.057297882e-07 wnfactor = -5.684341886e-20
+ eta0 = -4.522078841e-01 leta0 = 2.250651974e-07 weta0 = 3.330669074e-22 peta0 = -8.326672685e-29
+ etab = -1.886870119e-03 letab = 4.335647182e-10
+ u0 = 3.793238696e-02 lu0 = -7.159788098e-9
+ ua = 3.372214182e-09 lua = -1.059749752e-15 wua = -1.323488980e-29 pua = -3.308722450e-36
+ ub = 1.910230175e-18 lub = -4.885004854e-26
+ uc = -9.356751888e-11 luc = 2.211403977e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.213840779e+04 lvsat = 8.453340684e-3
+ a0 = 1.590800918e+00 la0 = -2.329470036e-7
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 2.018182291e-01 la2 = 1.419374407e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.486585336e-02 lketa = 5.541269763e-09 wketa = 4.440892099e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.369246124e-01 lpclm = 9.561406851e-8
+ pdiblc1 = -2.499817842e-01 lpdiblc1 = 1.563670691e-07 ppdiblc1 = -4.440892099e-28
+ pdiblc2 = -6.623202468e-03 lpdiblc2 = 3.630755750e-09 wpdiblc2 = -1.387778781e-23
+ pdiblcb = -1.647857919e-01 lpdiblcb = -2.943691991e-8
+ drout = 4.960126660e-01 ldrout = 7.803530650e-9
+ pscbe1 = -4.939454606e+08 lpscbe1 = 3.090783733e+02 ppscbe1 = -4.768371582e-19
+ pscbe2 = 1.444184156e-07 lpscbe2 = -3.238448899e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.995122502e+00 lbeta0 = 2.185239603e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.784636910e-09 lagidl = -4.259231038e-16
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.466034832e-01 lkt1 = -1.822337077e-8
+ kt2 = -6.597515796e-02 lkt2 = 3.144000191e-9
+ at = 9.157306403e+04 lat = -5.657723812e-3
+ ute = 3.308550878e-01 lute = -2.783895088e-7
+ ua1 = 2.975146297e-09 lua1 = -6.401978981e-16
+ ub1 = -1.532522831e-18 lub1 = 3.256279136e-25 pub1 = 3.081487911e-45
+ uc1 = -3.817149149e-11 luc1 = -1.426400859e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.160 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.367854064e-01 lvth0 = -4.651500081e-8
+ k1 = -6.134766510e-01 lk1 = 2.845755181e-7
+ k2 = 4.624846070e-01 lk2 = -1.135738648e-07 wk2 = -4.440892099e-22 pk2 = 1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.630409017e+00 ldsub = -2.020405853e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.162147361e-01 lvoff = -8.686492591e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.508360907e+00 lnfactor = 4.105193916e-7
+ eta0 = 4.900000007e-01 leta0 = -5.142197779e-17
+ etab = 1.809698392e-03 letab = -4.494346021e-10 wetab = -3.469446952e-24 petab = -4.336808690e-31
+ u0 = 1.773955312e-02 lu0 = -2.336325879e-9
+ ua = 1.258985607e-09 lua = -5.549628425e-16
+ ub = 8.412917613e-19 lub = 2.064872702e-25
+ uc = 2.878584554e-11 luc = -7.112508390e-18 wuc = 2.584939414e-32 puc = -3.231174268e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.331995797e+05 lvsat = -1.329844146e-2
+ a0 = -1.533380897e-02 la0 = 1.507103985e-7
+ ags = 2.122259360e+00 lags = -1.472984367e-7
+ a1 = 0.0
+ a2 = 9.101975611e-01 la2 = -2.727313031e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.777436513e-02 lketa = 1.101342597e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.768355118e-01 lpclm = -9.467448044e-9
+ pdiblc1 = 5.241829513e-01 lpdiblc1 = -2.855766128e-8
+ pdiblc2 = 2.628226065e-02 lpdiblc2 = -4.229372224e-9
+ pdiblcb = 1.765059758e+00 lpdiblcb = -4.904191263e-07 ppdiblcb = 8.881784197e-28
+ drout = -6.083418313e-01 ldrout = 2.716006894e-7
+ pscbe1 = 7.999088729e+08 lpscbe1 = 1.538864396e-2
+ pscbe2 = 1.774695567e-08 lpscbe2 = -2.126477355e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025125765e+01 lbeta0 = -3.203990428e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.492345636e-09 lagidl = 5.957197170e-16 wagidl = 2.791734567e-30 pagidl = -1.363555541e-36
+ bgidl = 1.818113540e+09 lbgidl = -1.381548262e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.689885319e-01 lkt1 = -3.676325419e-8
+ kt2 = -5.770354749e-02 lkt2 = 1.168160598e-9
+ at = 1.875627065e+05 lat = -2.858676971e-02 wat = 1.862645149e-15
+ ute = -1.682167421e+00 lute = 2.024611778e-7
+ ua1 = 1.624877580e-10 lua1 = 3.166184703e-17
+ ub1 = -3.030938486e-19 lub1 = 3.195421259e-26
+ uc1 = -2.633424711e-10 luc1 = 3.952258331e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.161 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 1.319595343e+01 lvth0 = -2.659462793e-06 wvth0 = -9.810007999e-06 pvth0 = 1.823386187e-12
+ k1 = 3.437067510e-01 lk1 = 1.353118157e-07 wk1 = 4.991269153e-07 pk1 = -9.277271974e-14
+ k2 = 1.055565439e+00 lk2 = -2.352431839e-07 wk2 = -8.677457269e-07 pk2 = 1.612878983e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.620398257e+00 ldsub = 9.394577079e-07 wdsub = 3.465394364e-06 pdsub = -6.441128505e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 3.579383892e+01 lvoff = -6.727009551e-06 wvoff = -2.481404066e-05 pvoff = 4.612185738e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -5.953739855e+02 lnfactor = 1.113943678e-04 wnfactor = 4.109024008e-04 pnfactor = -7.637442923e-11
+ eta0 = -9.842613315e+00 leta0 = 1.920522837e-06 weta0 = 7.084267008e-06 peta0 = -1.316752709e-12
+ etab = -5.875667322e-01 letab = 1.090527184e-07 wetab = 4.022646806e-07 petab = -7.476893618e-14
+ u0 = -6.007835564e-01 lu0 = 1.123933685e-07 wu0 = 4.145874231e-07 pu0 = -7.705936433e-14
+ ua = -1.174785227e-07 lua = 2.145891019e-14 wua = 7.915586642e-14 pua = -1.471270089e-20
+ ub = -4.918008739e-18 lub = 1.297755353e-24 wub = 4.787053471e-24 pub = -8.897696287e-31
+ uc = 4.392686841e-10 luc = -8.412496379e-17 wuc = -3.103132565e-16 puc = 5.767792498e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.284976480e+05 lvsat = -1.376323625e-02 wvsat = -5.076869469e-02 pvsat = 9.436377282e-9
+ a0 = 5.489747630e+00 la0 = -8.573472002e-07 wa0 = -3.162511241e-06 pa0 = 5.878159644e-13
+ ags = 1.250000057e+00 lags = -8.980734378e-15 wags = -2.601666438e-15 pags = 4.835811751e-22
+ a1 = 0.0
+ a2 = 7.800522124e+00 la2 = -1.310723320e-06 wa2 = -4.834888570e-06 pa2 = 8.986607385e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.804089990e+00 lketa = -3.376599895e-07 wketa = -1.245532441e-06 pketa = 2.315071148e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.592526162e-01 lpclm = -7.152395213e-09 wpclm = -2.638315620e-08 ppclm = 4.903837243e-15
+ pdiblc1 = -5.851099153e+00 lpdiblc1 = 1.153541148e-06 wpdiblc1 = 4.255088126e-06 ppdiblc1 = -7.908932300e-13
+ pdiblc2 = 3.108731910e-02 lpdiblc2 = -5.548255762e-09 wpdiblc2 = -2.046595435e-08 ppdiblc2 = 3.804006935e-15
+ pdiblcb = 3.493143043e+01 lpdiblcb = -6.704422521e-06 wpdiblcb = -2.473072352e-05 ppdiblcb = 4.596699581e-12
+ drout = 1.000000036e+00 ldrout = -1.875079647e-15 wdrout = 8.533254459e-14 pdrout = -1.586076337e-20
+ pscbe1 = 1.476796236e+08 lpscbe1 = 1.212467884e+02 wpscbe1 = 4.472452013e+02 ppscbe1 = -8.312946557e-5
+ pscbe2 = 1.417570559e-07 lpscbe2 = -2.539030536e-14 wpscbe2 = -9.365767662e-14 ppscbe2 = 1.740815235e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -3.902194178e+00 lbeta0 = 2.278048748e-06 wbeta0 = 8.403078730e-06 pbeta0 = -1.561880244e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.623997061e-07 lagidl = 6.755167141e-14 wagidl = 2.491790599e-13 pagidl = -4.631491186e-20
+ bgidl = 1.000000367e+09 lbgidl = -6.008681488e-05 wbgidl = -6.621429443e-05 pbgidl = 1.230725861e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.651281751e-02 lkt1 = -9.110924091e-08 wkt1 = -3.360764431e-07 pkt1 = 6.246652848e-14
+ kt2 = -1.487385738e+00 lkt2 = 2.670207870e-07 wkt2 = 9.849642433e-07 pkt2 = -1.830753039e-13
+ at = 1.288639548e+06 lat = -2.361217281e-01 wat = -8.709864303e-01 pat = 1.618902478e-7
+ ute = 1.036607634e+01 lute = -2.016564294e-06 wute = -7.438536998e-06 pute = 1.382600872e-12
+ ua1 = 1.369256582e-08 lua1 = -2.479986390e-15 wua1 = -9.147969564e-15 pua1 = 1.700333103e-21
+ ub1 = -1.819992810e-17 lub1 = 3.361655598e-24 wub1 = 1.240019885e-23 pub1 = -2.304824961e-30
+ uc1 = -4.392397940e-10 luc1 = 7.619532374e-17 wuc1 = 2.810630581e-16 puc1 = -5.224119061e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.162 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.163 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108623478e+00 lvth0 = 3.532668562e-7
+ k1 = 4.171052081e-01 lk1 = 2.908460917e-7
+ k2 = 2.159455618e-02 lk2 = -4.690448662e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 2.117582368e-27 pcit = 4.743384505e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.807199248e-01 lvoff = 2.151443021e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.403205388e+00 lnfactor = -5.131826301e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.149534990e-02 lu0 = -1.176644632e-8
+ ua = -9.044296180e-10 lua = 2.075453526e-15
+ ub = 1.700362603e-18 lub = -5.753769297e-24 wub = 1.540743956e-39
+ uc = -1.046578370e-10 luc = -2.009187197e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.286628951e+04 lvsat = -2.540643246e-1
+ a0 = 1.625827411e+00 la0 = -3.234747073e-6
+ ags = 1.127460711e-01 lags = 1.087252350e-8
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = -2.227955321e-07 lb0 = 2.397975426e-12 pb0 = -8.470329473e-34
+ b1 = 3.393294966e-09 lb1 = -2.149792907e-14
+ keta = 3.416681995e-02 lketa = -2.159909532e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 wpclm = -2.775557562e-23 ppclm = 6.661338148e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.906905271e-03 lpdiblc2 = -1.258792035e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.865952071e-09 lpscbe2 = 2.388016187e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.797495750e+01 lbeta0 = -3.592990887e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.808012713e-09 lagidl = -1.814500294e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443649873e-01 lkt1 = 1.222316870e-07 wkt1 = -4.440892099e-22
+ kt2 = -6.519461656e-02 lkt2 = 1.328983321e-7
+ at = 7.713361212e+04 lat = -1.228038641e-1
+ ute = 5.595779957e-01 lute = -1.284400824e-05 wute = -2.220446049e-22 pute = 4.440892099e-27
+ ua1 = 3.768264800e-09 lua1 = -3.354261913e-14
+ ub1 = -2.642787222e-18 lub1 = 2.826200788e-23 pub1 = 1.232595164e-44
+ uc1 = -9.417115820e-11 luc1 = 1.286926591e-15 wuc1 = -5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.164 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.068784975e+00 lvth0 = 3.500223376e-8
+ k1 = 4.603509166e-01 lk1 = -5.463825109e-8
+ k2 = 1.538364979e-02 lk2 = 2.713637080e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.682810246e-01 lvoff = 1.157715452e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.131821908e+00 lnfactor = 5.025091038e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.814547492e-03 lu0 = 9.650135606e-9
+ ua = -8.481377777e-10 lua = 1.625745332e-15
+ ub = 1.054996270e-18 lub = -5.980215607e-25
+ uc = -1.070085284e-10 luc = -1.312504100e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342054363e+04 lvsat = -1.882608877e-2
+ a0 = 1.169648264e+00 la0 = 4.096088288e-7
+ ags = 4.536500838e-02 lags = 5.491710742e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 5.989974384e-08 lb0 = 1.395596165e-13
+ b1 = -9.045963073e-10 lb1 = 1.283736559e-14 pb1 = 3.308722450e-36
+ keta = 7.536869066e-03 lketa = -3.247737421e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.061808156e-01 lpclm = 4.371028699e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.327209668e-04 lpdiblc2 = 7.869204170e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461096001e-08 lpscbe2 = -2.201595970e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.997217500e-10 lalpha0 = -7.966640969e-16
+ alpha1 = 1.997217500e-10 lalpha1 = -7.966640969e-16
+ beta0 = -2.392487250e+01 lbeta0 = 2.150993062e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.932747516e-10 lagidl = -1.250636281e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.139217330e-01 lkt1 = -1.209755144e-7
+ kt2 = -3.860015032e-02 lkt2 = -7.956140140e-8
+ at = 2.264263863e+04 lat = 3.125174394e-1
+ ute = -1.910932237e+00 lute = 6.892576840e-06 pute = 7.105427358e-27
+ ua1 = -2.943994399e-09 lua1 = 2.008074701e-14
+ ub1 = 2.913039917e-18 lub1 = -1.612277288e-23
+ uc1 = 5.506278879e-10 luc1 = -3.864289165e-15 wuc1 = -1.033975766e-31 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.165 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.063486545e+00 lvth0 = 1.386748510e-8
+ k1 = 3.863911154e-01 lk1 = 2.403777808e-7
+ k2 = 3.756574616e-02 lk2 = -8.576786165e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.583304901e-01 ldsub = -1.190001542e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.481840352e-01 lvoff = 3.560726699e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.206074825e+00 lnfactor = 7.400358035e-7
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391132325e-01 letab = 2.756836997e-7
+ u0 = 1.129796699e-02 lu0 = -2.559019068e-10
+ ua = -3.948101738e-10 lua = -1.825195469e-16
+ ub = 9.047694627e-19 lub = 1.213642946e-27
+ uc = -1.333555795e-10 luc = 1.037824576e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.345823238e+04 lvsat = -9.875382428e-2
+ a0 = 1.398566000e+00 la0 = -5.035142625e-7
+ ags = -4.042771799e-02 lags = 8.913871067e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 7.545275679e-08 lb0 = 7.752066969e-14
+ b1 = 6.234956092e-09 lb1 = -1.564138079e-14 pb1 = 6.617444900e-36
+ keta = 2.253544784e-02 lketa = -6.307511832e-08 wketa = -1.387778781e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.074223900e-01 lpclm = 3.278972801e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.187393462e-04 lpdiblc2 = 4.491728403e-11
+ pdiblcb = -4.238870000e-01 lpdiblcb = 7.933343877e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.718970657e-09 lpscbe2 = 1.486419869e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.944350000e-11 lalpha0 = 3.966671938e-16
+ alpha1 = -9.944350000e-11 lalpha1 = 3.966671938e-16
+ beta0 = 5.429614004e+01 lbeta0 = -9.691414411e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.573122120e-11 lagidl = 1.776939874e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356779703e-01 lkt1 = -3.419271211e-8
+ kt2 = -6.313133978e-02 lkt2 = 1.829032431e-8
+ at = 1.615988244e+05 lat = -2.417607213e-1
+ ute = -9.311290905e-02 lute = -3.584681431e-7
+ ua1 = 2.873317563e-09 lua1 = -3.123754152e-15
+ ub1 = -1.891532202e-18 lub1 = 3.042040710e-24
+ uc1 = -8.692813487e-10 luc1 = 1.799544192e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.166 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.081021165e+00 lvth0 = 4.874156567e-8
+ k1 = 5.064919019e-01 lk1 = 1.512929702e-9
+ k2 = -5.250837621e-03 lk2 = -6.112426770e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000199e-01 ldsub = -1.966733887e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.231624387e-01 lvoff = -1.415743548e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.405520147e+00 lnfactor = 3.433649873e-7
+ eta0 = -4.835518650e-01 leta0 = 9.627162327e-07 weta0 = -3.122502257e-23 peta0 = 3.747002708e-28
+ etab = 2.386594872e-04 letab = -1.469097694e-9
+ u0 = 1.277578903e-02 lu0 = -3.195097838e-9
+ ua = -2.787126111e-10 lua = -4.134225064e-16
+ ub = 8.338866336e-19 lub = 1.421903751e-25
+ uc = -1.183445084e-10 luc = 7.392738859e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.599790864e+04 lvsat = 3.541598979e-2
+ a0 = 1.034813481e+00 la0 = 2.199422095e-7
+ ags = 2.529917783e-01 lags = 3.078138731e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.221234086e-07 lb0 = -1.530118956e-14
+ b1 = -1.258163080e-08 lb1 = 2.178236438e-14 pb1 = 3.308722450e-36
+ keta = -1.722971284e-02 lketa = 1.601261680e-08 wketa = -1.387778781e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.149196182e-01 lpclm = -2.836747322e-07 wpclm = -8.881784197e-22
+ pdiblc1 = 3.955978546e-01 lpdiblc1 = -1.113340513e-8
+ pdiblc2 = 4.525213076e-04 lpdiblc2 = -2.227064540e-11
+ pdiblcb = 1.727740000e-01 lpdiblcb = -3.933467754e-07 ppdiblcb = -1.110223025e-28
+ drout = 3.855974777e-01 ldrout = 3.468639446e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.759262277e-09 lpscbe2 = -5.825849256e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.674544110e+00 lbeta0 = 1.776759381e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.258387184e-10 lagidl = 7.992711679e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.269668075e-01 lkt1 = -5.151808255e-8
+ kt2 = -5.925098613e-02 lkt2 = 1.057280534e-8
+ at = 2.845269774e+04 lat = 2.304961559e-2
+ ute = 4.928361669e-01 lute = -1.523844682e-6
+ ua1 = 3.016514543e-09 lua1 = -3.408554329e-15
+ ub1 = -1.565341614e-18 lub1 = 2.393290035e-24
+ uc1 = 4.482619664e-12 luc1 = 6.174124785e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.167 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.050737288e+00 lvth0 = 1.879474788e-8
+ k1 = 5.794701714e-01 lk1 = -7.065309168e-8
+ k2 = -3.599095491e-02 lk2 = 2.978673710e-08 wk2 = -6.938893904e-24 pk2 = 1.040834086e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.635276000e-01 ldsub = 7.154747378e-07 pdsub = -2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.308165965e-01 lvoff = -6.588468460e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.932418197e-01 lnfactor = 2.333246657e-6
+ eta0 = 9.611039418e-01 leta0 = -4.658605549e-7
+ etab = -1.488450021e-03 letab = 2.387890846e-10
+ u0 = -3.891442511e-03 lu0 = 1.328662742e-08 pu0 = -6.938893904e-30
+ ua = -2.555715282e-09 lua = 1.838237125e-15 wua = -8.271806126e-31 pua = 8.271806126e-37
+ ub = 1.635833473e-19 lub = 8.050331859e-25
+ uc = -3.894326448e-11 luc = -4.590119479e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.436459522e+04 lvsat = 7.365024437e-3
+ a0 = 1.396980751e+00 la0 = -1.381941390e-7
+ ags = -1.061952942e-01 lags = 6.630031935e-7
+ a1 = 0.0
+ a2 = 1.100991363e+00 la2 = -2.976413294e-07 wa2 = -8.881784197e-22
+ b0 = 2.109259710e-07 lb0 = -1.031153794e-13
+ b1 = 1.868153427e-08 lb1 = -9.132841657e-15
+ keta = 4.051134126e-02 lketa = -4.108577937e-08 wketa = 1.734723476e-24 pketa = 8.673617380e-30
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.192448538e-01 lpclm = -1.890648279e-7
+ pdiblc1 = 6.918059423e-01 lpdiblc1 = -3.040446968e-07 wpdiblc1 = -4.440892099e-22
+ pdiblc2 = 6.468668115e-05 lpdiblc2 = 3.612473816e-10
+ pdiblcb = -0.225
+ drout = 9.557609593e-01 ldrout = -2.169536175e-07 wdrout = -8.881784197e-22
+ pscbe1 = 1.446985488e+09 lpscbe1 = -6.397845396e+02 ppscbe1 = 4.768371582e-19
+ pscbe2 = -5.829857018e-08 lpscbe2 = 6.671776386e-14 ppscbe2 = -2.646977960e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.544352635e+00 lbeta0 = 1.905501825e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.547675918e-09 lagidl = -3.100799834e-16 wagidl = -1.654361225e-30
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.743566677e-01 lkt1 = -4.655671468e-9
+ kt2 = -3.781888407e-02 lkt2 = -1.062075742e-8
+ at = 2.415206960e+04 lat = 2.730237773e-2
+ ute = -1.839698799e+00 lute = 7.827291698e-7
+ ua1 = -2.479750931e-09 lua1 = 2.026537710e-15 pua1 = -4.135903063e-37
+ ub1 = 2.537894393e-18 lub1 = -1.664276955e-24
+ uc1 = 1.981977632e-10 luc1 = -1.298178461e-16 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.168 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.939250368e-01 lvth0 = -8.979057300e-9
+ k1 = 2.983925622e-01 lk1 = 6.675731910e-8
+ k2 = 6.116802299e-02 lk2 = -1.771137242e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.205819134e+00 ldsub = -1.006188000e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.412922644e-01 lvoff = -1.467228692e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.018676894e+00 lnfactor = -9.057297882e-07 wnfactor = -7.105427358e-21
+ eta0 = -4.522078841e-01 leta0 = 2.250651974e-07 weta0 = -1.526556659e-22 peta0 = -5.204170428e-29
+ etab = -1.886870119e-03 letab = 4.335647182e-10
+ u0 = 3.793238696e-02 lu0 = -7.159788098e-9
+ ua = 3.372214182e-09 lua = -1.059749752e-15 pua = -4.135903063e-37
+ ub = 1.910230175e-18 lub = -4.885004854e-26
+ uc = -9.356751888e-11 luc = 2.211403977e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.213840779e+04 lvsat = 8.453340684e-3
+ a0 = 1.590800918e+00 la0 = -2.329470036e-7
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 2.018182291e-01 la2 = 1.419374407e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.486585336e-02 lketa = 5.541269763e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.369246124e-01 lpclm = 9.561406851e-8
+ pdiblc1 = -2.499817842e-01 lpdiblc1 = 1.563670691e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = 5.551115123e-29
+ pdiblc2 = -6.623202468e-03 lpdiblc2 = 3.630755750e-09 wpdiblc2 = -1.734723476e-24 ppdiblc2 = -6.505213035e-31
+ pdiblcb = -1.647857919e-01 lpdiblcb = -2.943691991e-8
+ drout = 4.960126660e-01 ldrout = 7.803530650e-9
+ pscbe1 = -4.939454606e+08 lpscbe1 = 3.090783733e+02 ppscbe1 = 5.960464478e-20
+ pscbe2 = 1.444184156e-07 lpscbe2 = -3.238448899e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.995122502e+00 lbeta0 = 2.185239603e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.784636910e-09 lagidl = -4.259231038e-16
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.466034832e-01 lkt1 = -1.822337077e-8
+ kt2 = -6.597515796e-02 lkt2 = 3.144000191e-9
+ at = 9.157306403e+04 lat = -5.657723812e-3
+ ute = 3.308550878e-01 lute = -2.783895088e-07 pute = 1.110223025e-28
+ ua1 = 2.975146297e-09 lua1 = -6.401978981e-16
+ ub1 = -1.532522831e-18 lub1 = 3.256279136e-25
+ uc1 = -3.817149149e-11 luc1 = -1.426400859e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.169 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.367854064e-01 lvth0 = -4.651500081e-8
+ k1 = -6.134766510e-01 lk1 = 2.845755181e-7
+ k2 = 4.624846070e-01 lk2 = -1.135738648e-07 wk2 = 5.551115123e-23 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.630409017e+00 ldsub = -2.020405853e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.162147361e-01 lvoff = -8.686492591e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.508360907e+00 lnfactor = 4.105193916e-7
+ eta0 = 4.900000007e-01 leta0 = -5.142020143e-17
+ etab = 1.809698392e-03 letab = -4.494346021e-10 wetab = 8.673617380e-25 petab = 1.355252716e-31
+ u0 = 1.773955312e-02 lu0 = -2.336325879e-9
+ ua = 1.258985607e-09 lua = -5.549628425e-16
+ ub = 8.412917613e-19 lub = 2.064872702e-25
+ uc = 2.878584554e-11 luc = -7.112508390e-18 wuc = 9.693522803e-33 puc = -1.615587134e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.331995797e+05 lvsat = -1.329844146e-2
+ a0 = -1.533380897e-02 la0 = 1.507103985e-7
+ ags = 2.122259360e+00 lags = -1.472984367e-7
+ a1 = 0.0
+ a2 = 9.101975611e-01 la2 = -2.727313031e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.777436513e-02 lketa = 1.101342597e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.768355118e-01 lpclm = -9.467448044e-9
+ pdiblc1 = 5.241829513e-01 lpdiblc1 = -2.855766128e-8
+ pdiblc2 = 2.628226065e-02 lpdiblc2 = -4.229372224e-9
+ pdiblcb = 1.765059758e+00 lpdiblcb = -4.904191263e-07 wpdiblcb = -8.881784197e-22
+ drout = -6.083418313e-01 ldrout = 2.716006894e-7
+ pscbe1 = 7.999088729e+08 lpscbe1 = 1.538864396e-2
+ pscbe2 = 1.774695567e-08 lpscbe2 = -2.126477355e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025125765e+01 lbeta0 = -3.203990428e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.492345636e-09 lagidl = 5.957197170e-16 wagidl = -6.009984138e-31 pagidl = -1.866003140e-37
+ bgidl = 1.818113540e+09 lbgidl = -1.381548262e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.689885319e-01 lkt1 = -3.676325419e-8
+ kt2 = -5.770354749e-02 lkt2 = 1.168160598e-9
+ at = 1.875627065e+05 lat = -2.858676971e-02 pat = 2.910383046e-23
+ ute = -1.682167421e+00 lute = 2.024611778e-7
+ ua1 = 1.624877580e-10 lua1 = 3.166184703e-17
+ ub1 = -3.030938486e-19 lub1 = 3.195421259e-26
+ uc1 = -2.633424711e-10 luc1 = 3.952258331e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.170 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -2.395090936e+00 lvth0 = 2.384446222e-07 wvth0 = 7.236445746e-07 pvth0 = -1.345038171e-13
+ k1 = 3.319605812e-01 lk1 = 1.374950763e-07 wk1 = 5.070628860e-07 pk1 = -9.424777862e-14
+ k2 = -1.793692352e-01 lk2 = -5.705876060e-09 wk2 = -3.339669248e-08 pk2 = 6.207443231e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.701950988e+00 ldsub = 9.546159140e-07 wdsub = 3.520493183e-06 pdsub = -6.543540680e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -4.550210120e+00 lvoff = 7.717388435e-07 wvoff = 2.443286439e-06 pvoff = -4.541336504e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.233373617e+01 lnfactor = -1.271246647e-05 wnfactor = -4.021562561e-05 pnfactor = 7.474878332e-12
+ eta0 = -1.000933158e+01 leta0 = 1.951510761e-06 weta0 = 7.196905538e-06 peta0 = -1.337688832e-12
+ etab = -5.970333503e-01 letab = 1.108122787e-07 wetab = 4.086605360e-07 petab = -7.595773382e-14
+ u0 = 7.270932895e-02 lu0 = -1.278875406e-08 wu0 = -4.043918710e-08 pu0 = 7.516431706e-15
+ ua = 8.588555829e-09 lua = -1.973177699e-15 wua = -6.017825308e-15 pua = 1.118533190e-21
+ ub = 7.278130866e-18 lub = -9.691411154e-25 wub = -3.452926761e-24 pub = 6.417954971e-31
+ uc = 4.465714238e-10 luc = -8.548232402e-17 wuc = -3.152471481e-16 puc = 5.859498742e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.339396742e+05 lvsat = 7.218998882e-02 wvsat = 2.616641338e-01 pvsat = -4.863551255e-8
+ a0 = 5.564172799e+00 la0 = -8.711806064e-07 wa0 = -3.212794523e-06 pa0 = 5.971621179e-13
+ ags = 1.250000053e+00 lags = -8.187253542e-15 wags = 2.825188972e-16 pags = -5.251177271e-23
+ a1 = 0.0
+ a2 = 7.914304040e+00 la2 = -1.331871965e-06 wa2 = -4.911762136e-06 pa2 = 9.129492282e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.833401555e+00 lketa = -3.431081300e-07 wketa = -1.265335979e-06 pketa = 2.351879984e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.598735084e-01 lpclm = -7.267800440e-09 wpclm = -2.680264461e-08 ppclm = 4.981807553e-15
+ pdiblc1 = -5.951236129e+00 lpdiblc1 = 1.172153608e-06 wpdiblc1 = 4.322742870e-06 ppdiblc1 = -8.034682172e-13
+ pdiblc2 = 3.156894820e-02 lpdiblc2 = -5.637776163e-09 wpdiblc2 = -2.079135357e-08 ppdiblc2 = 3.864488888e-15
+ pdiblcb = 3.551343339e+01 lpdiblcb = -6.812599412e-06 wpdiblcb = -2.512393753e-05 ppdiblcb = 4.669786268e-12
+ drout = 1.000000176e+00 ldrout = -2.790014442e-14 wdrout = -9.266393874e-15 pdrout = 1.722344045e-21
+ pscbe1 = 1.371544465e+08 lpscbe1 = 1.232031030e+02 wpscbe1 = 4.543562426e+02 ppscbe1 = -8.445119480e-5
+ pscbe2 = 1.439611197e-07 lpscbe2 = -2.579997469e-14 wpscbe2 = -9.514679060e-14 ppscbe2 = 1.768493397e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -4.099948165e+00 lbeta0 = 2.314805282e-06 wbeta0 = 8.536685675e-06 pbeta0 = -1.586713766e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.780010855e-08 lagidl = -8.692168143e-15 wagidl = -2.796095931e-14 pagidl = 5.197103506e-21
+ bgidl = 1.000000258e+09 lbgidl = -3.989249611e-05 wbgidl = 7.190319061e-06 pbgidl = -1.336463928e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.860385105e-02 lkt1 = -9.257928051e-08 wkt1 = -3.414199148e-07 pkt1 = 6.345971957e-14
+ kt2 = -1.510565206e+00 lkt2 = 2.713291548e-07 wkt2 = 1.000624802e-06 pkt2 = -1.859861320e-13
+ at = 1.309136784e+06 lat = -2.399315494e-01 wat = -8.848348139e-01 pat = 1.644642469e-7
+ ute = 1.054113156e+01 lute = -2.049101809e-06 wute = -7.556808160e-06 pute = 1.404583933e-12
+ ua1 = 1.390785269e-08 lua1 = -2.520001761e-15 wua1 = -9.293422110e-15 pua1 = 1.727368368e-21
+ ub1 = -1.849174368e-17 lub1 = 3.415895360e-24 wub1 = 1.259735588e-23 pub1 = -2.341470537e-30
+ uc1 = -4.458541873e-10 luc1 = 7.742474102e-17 wuc1 = 2.855318877e-16 puc1 = -5.307181197e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.171 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.172 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.108623478e+00 lvth0 = 3.532668562e-07 wvth0 = 7.105427358e-21
+ k1 = 4.171052081e-01 lk1 = 2.908460917e-7
+ k2 = 2.159455618e-02 lk2 = -4.690448662e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 1.355252716e-26 pcit = 1.084202172e-31
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.807199248e-01 lvoff = 2.151443021e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.403205388e+00 lnfactor = -5.131826301e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.149534990e-02 lu0 = -1.176644632e-8
+ ua = -9.044296180e-10 lua = 2.075453526e-15
+ ub = 1.700362603e-18 lub = -5.753769297e-24
+ uc = -1.046578370e-10 luc = -2.009187197e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.286628951e+04 lvsat = -2.540643246e-1
+ a0 = 1.625827411e+00 la0 = -3.234747073e-6
+ ags = 1.127460711e-01 lags = 1.087252350e-8
+ a1 = 0.0
+ a2 = 1.083175658e+00 la2 = -2.262253522e-6
+ b0 = -2.227955321e-07 lb0 = 2.397975426e-12 pb0 = -6.776263578e-33
+ b1 = 3.393294966e-09 lb1 = -2.149792907e-14
+ keta = 3.416681995e-02 lketa = -2.159909532e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.885582638e-02 lpclm = 1.676183212e-06 wpclm = -1.110223025e-22 ppclm = 3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.906905271e-03 lpdiblc2 = -1.258792035e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.865952071e-09 lpscbe2 = 2.388016187e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.657391667e-11 lalpha0 = 1.330737366e-15
+ alpha1 = -6.657391667e-11 lalpha1 = 1.330737366e-15
+ beta0 = 4.797495750e+01 lbeta0 = -3.592990887e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.808012713e-09 lagidl = -1.814500294e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443649873e-01 lkt1 = 1.222316870e-7
+ kt2 = -6.519461656e-02 lkt2 = 1.328983321e-7
+ at = 7.713361212e+04 lat = -1.228038641e-1
+ ute = 5.595779957e-01 lute = -1.284400824e-05 pute = -1.421085472e-26
+ ua1 = 3.768264800e-09 lua1 = -3.354261913e-14
+ ub1 = -2.642787222e-18 lub1 = 2.826200788e-23 pub1 = 9.860761315e-44
+ uc1 = -9.417115820e-11 luc1 = 1.286926591e-15 puc1 = 3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.173 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.068784975e+00 lvth0 = 3.500223376e-8
+ k1 = 4.603509166e-01 lk1 = -5.463825109e-8
+ k2 = 1.538364979e-02 lk2 = 2.713637080e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.682810246e-01 lvoff = 1.157715452e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.131821908e+00 lnfactor = 5.025091038e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.814547492e-03 lu0 = 9.650135606e-9
+ ua = -8.481377777e-10 lua = 1.625745332e-15
+ ub = 1.054996270e-18 lub = -5.980215607e-25
+ uc = -1.070085284e-10 luc = -1.312504100e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342054363e+04 lvsat = -1.882608877e-2
+ a0 = 1.169648264e+00 la0 = 4.096088288e-7
+ ags = 4.536500838e-02 lags = 5.491710742e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 5.989974383e-08 lb0 = 1.395596165e-13
+ b1 = -9.045963073e-10 lb1 = 1.283736559e-14 pb1 = 2.646977960e-35
+ keta = 7.536869066e-03 lketa = -3.247737421e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.061808156e-01 lpclm = 4.371028699e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.327209668e-04 lpdiblc2 = 7.869204170e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461096001e-08 lpscbe2 = -2.201595970e-14 wpscbe2 = -1.058791184e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.997217500e-10 lalpha0 = -7.966640969e-16
+ alpha1 = 1.997217500e-10 lalpha1 = -7.966640969e-16
+ beta0 = -2.392487250e+01 lbeta0 = 2.150993062e-04 wbeta0 = 2.842170943e-20 pbeta0 = -3.410605132e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.932747516e-10 lagidl = -1.250636281e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.139217330e-01 lkt1 = -1.209755144e-7
+ kt2 = -3.860015032e-02 lkt2 = -7.956140140e-8
+ at = 2.264263863e+04 lat = 3.125174394e-1
+ ute = -1.910932237e+00 lute = 6.892576840e-6
+ ua1 = -2.943994399e-09 lua1 = 2.008074701e-14 wua1 = -6.617444900e-30 pua1 = 2.646977960e-35
+ ub1 = 2.913039917e-18 lub1 = -1.612277288e-23
+ uc1 = 5.506278879e-10 luc1 = -3.864289165e-15 wuc1 = -1.654361225e-30 puc1 = 9.926167351e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.174 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.063486545e+00 lvth0 = 1.386748510e-8
+ k1 = 3.863911154e-01 lk1 = 2.403777808e-7
+ k2 = 3.756574616e-02 lk2 = -8.576786165e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.583304901e-01 ldsub = -1.190001542e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.481840352e-01 lvoff = 3.560726699e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.206074825e+00 lnfactor = 7.400358035e-7
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391132325e-01 letab = 2.756836997e-7
+ u0 = 1.129796699e-02 lu0 = -2.559019068e-10
+ ua = -3.948101738e-10 lua = -1.825195469e-16
+ ub = 9.047694627e-19 lub = 1.213642946e-27
+ uc = -1.333555795e-10 luc = 1.037824576e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.345823238e+04 lvsat = -9.875382428e-2
+ a0 = 1.398566000e+00 la0 = -5.035142625e-7
+ ags = -4.042771799e-02 lags = 8.913871067e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 7.545275679e-08 lb0 = 7.752066969e-14
+ b1 = 6.234956092e-09 lb1 = -1.564138079e-14
+ keta = 2.253544784e-02 lketa = -6.307511832e-08 wketa = 5.551115123e-23 pketa = 1.110223025e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.074223900e-01 lpclm = 3.278972801e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.187393462e-04 lpdiblc2 = 4.491728403e-11
+ pdiblcb = -4.238870000e-01 lpdiblcb = 7.933343877e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.718970657e-09 lpscbe2 = 1.486419869e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.944350000e-11 lalpha0 = 3.966671938e-16
+ alpha1 = -9.944350000e-11 lalpha1 = 3.966671938e-16
+ beta0 = 5.429614004e+01 lbeta0 = -9.691414411e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.573122120e-11 lagidl = 1.776939874e-15 pagidl = 6.617444900e-36
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356779703e-01 lkt1 = -3.419271211e-8
+ kt2 = -6.313133979e-02 lkt2 = 1.829032431e-8
+ at = 1.615988244e+05 lat = -2.417607213e-1
+ ute = -9.311290905e-02 lute = -3.584681431e-7
+ ua1 = 2.873317562e-09 lua1 = -3.123754152e-15
+ ub1 = -1.891532202e-18 lub1 = 3.042040710e-24
+ uc1 = -8.692813487e-10 luc1 = 1.799544192e-15 puc1 = 6.617444900e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.175 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.081021165e+00 lvth0 = 4.874156567e-8
+ k1 = 5.064919019e-01 lk1 = 1.512929702e-9
+ k2 = -5.250837621e-03 lk2 = -6.112426770e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000199e-01 ldsub = -1.966733620e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.231624387e-01 lvoff = -1.415743548e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.405520147e+00 lnfactor = 3.433649873e-7
+ eta0 = -4.835518650e-01 leta0 = 9.627162327e-07 weta0 = -8.118505868e-22 peta0 = 2.851885395e-27
+ etab = 2.386594872e-04 letab = -1.469097694e-9
+ u0 = 1.277578903e-02 lu0 = -3.195097838e-9
+ ua = -2.787126111e-10 lua = -4.134225064e-16
+ ub = 8.338866336e-19 lub = 1.421903751e-25
+ uc = -1.183445084e-10 luc = 7.392738859e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.599790864e+04 lvsat = 3.541598979e-2
+ a0 = 1.034813481e+00 la0 = 2.199422095e-7
+ ags = 2.529917783e-01 lags = 3.078138731e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.221234086e-07 lb0 = -1.530118956e-14
+ b1 = -1.258163080e-08 lb1 = 2.178236438e-14 pb1 = 3.970466940e-35
+ keta = -1.722971284e-02 lketa = 1.601261680e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.149196182e-01 lpclm = -2.836747322e-7
+ pdiblc1 = 3.955978546e-01 lpdiblc1 = -1.113340513e-8
+ pdiblc2 = 4.525213076e-04 lpdiblc2 = -2.227064540e-11
+ pdiblcb = 1.727740000e-01 lpdiblcb = -3.933467754e-07 wpdiblcb = -2.220446049e-22 ppdiblcb = -4.440892099e-28
+ drout = 3.855974777e-01 ldrout = 3.468639446e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.759262277e-09 lpscbe2 = -5.825849256e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.674544110e+00 lbeta0 = 1.776759381e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.258387184e-10 lagidl = 7.992711679e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.269668075e-01 lkt1 = -5.151808255e-8
+ kt2 = -5.925098613e-02 lkt2 = 1.057280534e-8
+ at = 2.845269774e+04 lat = 2.304961559e-2
+ ute = 4.928361669e-01 lute = -1.523844682e-6
+ ua1 = 3.016514543e-09 lua1 = -3.408554329e-15
+ ub1 = -1.565341614e-18 lub1 = 2.393290035e-24 wub1 = -3.081487911e-39
+ uc1 = 4.482619664e-12 luc1 = 6.174124785e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.176 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.050737288e+00 lvth0 = 1.879474788e-8
+ k1 = 5.794701714e-01 lk1 = -7.065309168e-8
+ k2 = -3.599095491e-02 lk2 = 2.978673710e-08 wk2 = -5.551115123e-23 pk2 = 8.326672685e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.635276000e-01 ldsub = 7.154747378e-07 pdsub = -1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.308165965e-01 lvoff = -6.588468460e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.932418197e-01 lnfactor = 2.333246657e-6
+ eta0 = 9.611039418e-01 leta0 = -4.658605549e-7
+ etab = -1.488450021e-03 letab = 2.387890846e-10
+ u0 = -3.891442511e-03 lu0 = 1.328662742e-8
+ ua = -2.555715282e-09 lua = 1.838237125e-15 wua = 6.617444900e-30 pua = 3.308722450e-36
+ ub = 1.635833473e-19 lub = 8.050331859e-25
+ uc = -3.894326448e-11 luc = -4.590119479e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.436459522e+04 lvsat = 7.365024437e-3
+ a0 = 1.396980751e+00 la0 = -1.381941390e-7
+ ags = -1.061952942e-01 lags = 6.630031935e-7
+ a1 = 0.0
+ a2 = 1.100991363e+00 la2 = -2.976413294e-7
+ b0 = 2.109259710e-07 lb0 = -1.031153794e-13
+ b1 = 1.868153427e-08 lb1 = -9.132841657e-15
+ keta = 4.051134126e-02 lketa = -4.108577937e-08 wketa = 9.714451465e-23 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.192448538e-01 lpclm = -1.890648279e-7
+ pdiblc1 = 6.918059423e-01 lpdiblc1 = -3.040446968e-7
+ pdiblc2 = 6.468668115e-05 lpdiblc2 = 3.612473816e-10
+ pdiblcb = -0.225
+ drout = 9.557609593e-01 ldrout = -2.169536175e-7
+ pscbe1 = 1.446985488e+09 lpscbe1 = -6.397845396e+2
+ pscbe2 = -5.829857018e-08 lpscbe2 = 6.671776386e-14 wpscbe2 = -1.058791184e-28 ppscbe2 = -2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.544352635e+00 lbeta0 = 1.905501825e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.547675918e-09 lagidl = -3.100799834e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.743566677e-01 lkt1 = -4.655671468e-9
+ kt2 = -3.781888407e-02 lkt2 = -1.062075742e-8
+ at = 2.415206960e+04 lat = 2.730237773e-2
+ ute = -1.839698799e+00 lute = 7.827291698e-7
+ ua1 = -2.479750931e-09 lua1 = 2.026537710e-15 pua1 = -1.654361225e-36
+ ub1 = 2.537894393e-18 lub1 = -1.664276955e-24
+ uc1 = 1.981977632e-10 luc1 = -1.298178461e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.177 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.939250368e-01 lvth0 = -8.979057300e-9
+ k1 = 2.983925622e-01 lk1 = 6.675731910e-8
+ k2 = 6.116802299e-02 lk2 = -1.771137242e-08 wk2 = 2.220446049e-22
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.205819134e+00 ldsub = -1.006188000e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.412922644e-01 lvoff = -1.467228692e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 7.018676894e+00 lnfactor = -9.057297882e-7
+ eta0 = -4.522078841e-01 leta0 = 2.250651974e-07 weta0 = -7.771561172e-22 peta0 = 8.326672685e-29
+ etab = -1.886870119e-03 letab = 4.335647182e-10
+ u0 = 3.793238696e-02 lu0 = -7.159788098e-9
+ ua = 3.372214182e-09 lua = -1.059749752e-15 wua = -1.323488980e-29
+ ub = 1.910230175e-18 lub = -4.885004854e-26
+ uc = -9.356751888e-11 luc = 2.211403977e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.213840779e+04 lvsat = 8.453340684e-3
+ a0 = 1.590800918e+00 la0 = -2.329470036e-7
+ ags = 1.005767373e+00 lags = 1.193980042e-7
+ a1 = 0.0
+ a2 = 2.018182291e-01 la2 = 1.419374407e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.486585336e-02 lketa = 5.541269763e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.369246124e-01 lpclm = 9.561406851e-8
+ pdiblc1 = -2.499817842e-01 lpdiblc1 = 1.563670691e-07 wpdiblc1 = 8.881784197e-22 ppdiblc1 = -2.220446049e-28
+ pdiblc2 = -6.623202468e-03 lpdiblc2 = 3.630755750e-09 wpdiblc2 = -6.938893904e-24 ppdiblc2 = -1.040834086e-29
+ pdiblcb = -1.647857919e-01 lpdiblcb = -2.943691991e-8
+ drout = 4.960126660e-01 ldrout = 7.803530650e-9
+ pscbe1 = -4.939454606e+08 lpscbe1 = 3.090783733e+02 wpscbe1 = -1.907348633e-12 ppscbe1 = 9.536743164e-19
+ pscbe2 = 1.444184156e-07 lpscbe2 = -3.238448899e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.995122502e+00 lbeta0 = 2.185239603e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.784636910e-09 lagidl = -4.259231038e-16
+ bgidl = 7.709281792e+08 lbgidl = 1.119863410e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.466034832e-01 lkt1 = -1.822337077e-8
+ kt2 = -6.597515796e-02 lkt2 = 3.144000191e-9
+ at = 9.157306403e+04 lat = -5.657723812e-3
+ ute = 3.308550878e-01 lute = -2.783895088e-07 pute = -4.440892099e-28
+ ua1 = 2.975146297e-09 lua1 = -6.401978981e-16
+ ub1 = -1.532522831e-18 lub1 = 3.256279136e-25
+ uc1 = -3.817149149e-11 luc1 = -1.426400859e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.178 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -8.367854064e-01 lvth0 = -4.651500081e-8
+ k1 = -6.134766510e-01 lk1 = 2.845755181e-7
+ k2 = 4.624846070e-01 lk2 = -1.135738648e-07 wk2 = 8.881784197e-22 pk2 = 5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.630409017e+00 ldsub = -2.020405853e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 1.162147361e-01 lvoff = -8.686492591e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.508360907e+00 lnfactor = 4.105193916e-7
+ eta0 = 4.900000007e-01 leta0 = -5.141842507e-17
+ etab = 1.809698392e-03 letab = -4.494346021e-10 wetab = -5.204170428e-24 petab = -1.084202172e-30
+ u0 = 1.773955312e-02 lu0 = -2.336325879e-9
+ ua = 1.258985607e-09 lua = -5.549628425e-16
+ ub = 8.412917613e-19 lub = 2.064872702e-25
+ uc = 2.878584554e-11 luc = -7.112508390e-18 wuc = -5.169878828e-32 puc = -1.615587134e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.331995797e+05 lvsat = -1.329844146e-2
+ a0 = -1.533380897e-02 la0 = 1.507103985e-7
+ ags = 2.122259360e+00 lags = -1.472984367e-7
+ a1 = 0.0
+ a2 = 9.101975611e-01 la2 = -2.727313031e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.777436513e-02 lketa = 1.101342597e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.768355118e-01 lpclm = -9.467448044e-9
+ pdiblc1 = 5.241829513e-01 lpdiblc1 = -2.855766128e-8
+ pdiblc2 = 2.628226065e-02 lpdiblc2 = -4.229372224e-9
+ pdiblcb = 1.765059758e+00 lpdiblcb = -4.904191263e-07 ppdiblcb = 8.881784197e-28
+ drout = -6.083418313e-01 ldrout = 2.716006894e-7
+ pscbe1 = 7.999088729e+08 lpscbe1 = 1.538864396e-2
+ pscbe2 = 1.774695567e-08 lpscbe2 = -2.126477355e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.025125765e+01 lbeta0 = -3.203990428e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.492345636e-09 lagidl = 5.957197170e-16 wagidl = 1.757758802e-30 pagidl = -1.156760388e-36
+ bgidl = 1.818113540e+09 lbgidl = -1.381548262e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644019647032
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.29936672419988e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.689885319e-01 lkt1 = -3.676325419e-8
+ kt2 = -5.770354749e-02 lkt2 = 1.168160598e-9
+ at = 1.875627065e+05 lat = -2.858676971e-2
+ ute = -1.682167421e+00 lute = 2.024611778e-7
+ ua1 = 1.624877580e-10 lua1 = 3.166184703e-17
+ ub1 = -3.030938486e-19 lub1 = 3.195421259e-26
+ uc1 = -2.633424711e-10 luc1 = 3.952258331e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.179 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 9.725373491e+00 lvth0 = -2.014386101e-06 wvth0 = -6.495570688e-06 pvth0 = 1.207331724e-12
+ k1 = -2.258766977e-01 lk1 = 2.411802913e-07 wk1 = 8.393230418e-07 pk1 = -1.560049738e-13
+ k2 = -1.686043594e+00 lk2 = 2.743396871e-07 wk2 = 8.640117026e-07 pk2 = -1.605938552e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.848290830e+00 ldsub = -8.204875327e-07 wdsub = -2.167840949e-06 pdsub = 4.029365972e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 2.776934175e+01 lvoff = -5.235496263e-06 wvoff = -1.680694968e-05 pvoff = 3.123907738e-12
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -4.193396401e+02 lnfactor = 7.867486398e-05 wnfactor = 2.526358541e-04 pnfactor = -4.695742620e-11
+ eta0 = 7.565480815e+00 leta0 = -1.315119619e-06 weta0 = -3.271039372e-06 peta0 = 6.079880881e-13
+ etab = 4.049986945e-01 letab = -7.543541751e-08 wetab = -1.881717946e-07 petab = 3.497549146e-14
+ u0 = -3.180683585e-01 lu0 = 5.984509470e-08 wu0 = 1.923166006e-07 pu0 = -3.574588656e-14
+ ua = -1.891914974e-08 lua = 3.139679534e-15 wua = 1.036636930e-14 pua = -1.926797061e-21
+ ub = -5.744425811e-17 lub = 1.106080932e-23 wub = 3.509715201e-23 pub = -6.523507643e-30
+ uc = -4.282788327e-10 luc = 7.712609314e-17 wuc = 2.058329114e-16 puc = -3.825816323e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.016476799e+06 lvsat = -7.364219211e-01 wvsat = -2.329539627e+00 pvsat = 4.329915304e-7
+ a0 = 2.201214274e-02 la0 = 1.589407948e-07 wa0 = 8.823829167e-08 pa0 = -1.640085127e-14
+ ags = 1.249999926e+00 lags = 1.538647609e-14 wags = 7.582468697e-14 pags = -1.409353700e-20
+ a1 = 0.0
+ a2 = -6.144436002e+00 la2 = 1.281226047e-06 wa2 = 3.461932726e-06 pa2 = -6.434694357e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.340882724e+00 lketa = 2.468960890e-07 wketa = 6.253375723e-07 pketa = -1.162314946e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.628759095e-01 lpclm = -7.825856746e-09 wpclm = -2.859094080e-08 ppclm = 5.314198166e-15
+ pdiblc1 = 1.148677440e+00 lpdiblc1 = -1.475073275e-07 wpdiblc1 = 9.387815034e-08 ppdiblc1 = -1.744913180e-14
+ pdiblc2 = 2.527577101e-02 lpdiblc2 = -4.468063319e-09 wpdiblc2 = -1.704299878e-08 ppdiblc2 = 3.167782184e-15
+ pdiblcb = -1.443754083e+01 lpdiblcb = 2.471788166e-06 wpdiblcb = 4.627961642e-06 ppdiblcb = -8.601992303e-13
+ drout = 1.000000030e+00 ldrout = -8.456240153e-16 wdrout = 7.743003039e-14 pdrout = -1.439192232e-20
+ pscbe1 = 1.246682778e+09 lpscbe1 = -8.302492798e+01 wpscbe1 = -2.065032415e+02 ppscbe1 = 3.838275749e-5
+ pscbe2 = -1.060382373e-08 lpscbe2 = 2.929011338e-15 wpscbe2 = -3.084509878e-15 ppscbe2 = 5.733178510e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.725114145e+01 lbeta0 = -1.653721745e-06 wbeta0 = -4.180493024e-06 pbeta0 = 7.770282384e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.246694584e-07 lagidl = 6.053875026e-14 wagidl = 1.938901091e-13 pagidl = -3.603835458e-20
+ bgidl = 1.000000359e+09 lbgidl = -5.860388184e-05 wbgidl = -5.277047729e-05 pbgidl = 9.808448792e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.406670741e-01 lkt1 = -1.537808674e-07 wkt1 = -5.375409218e-07 pkt1 = 9.991273114e-14
+ kt2 = 9.691529664e-01 lkt2 = -1.895760619e-07 wkt2 = -4.763498952e-07 pkt2 = 8.853915502e-14
+ at = -5.116395771e+05 lat = 9.849615283e-02 wat = 1.996596437e-01 pat = -3.711073798e-8
+ ute = -2.146123259e+00 lute = 3.090782449e-07 wute = -6.872357972e-14 pute = 1.277365058e-20
+ ua1 = 1.104806946e-10 lua1 = 4.451577126e-17 wua1 = -1.075403810e-15 pua1 = 1.998853061e-22
+ ub1 = 2.980863316e-18 lub1 = -5.752181021e-25 wub1 = -1.922012433e-25 pub1 = 3.572444508e-32
+ uc1 = -7.122960440e-10 luc1 = 1.269482889e-16 wuc1 = 4.442305192e-16 puc1 = -8.256912661e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.180 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.181 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.142549029e+00 lvth0 = 1.031400288e-06 wvth0 = 1.986754912e-08 pvth0 = -3.971298566e-13
+ k1 = 3.602134186e-01 lk1 = 1.428048676e-06 wk1 = 3.331708355e-08 pk1 = -6.659708518e-13
+ k2 = 2.591525663e-02 lk2 = -1.332704063e-07 wk2 = -2.530297242e-09 pk2 = 5.057778264e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = 6.352747104e-28 pcit = -1.863472484e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -3.087347497e-01 lvoff = 7.751289954e-07 wvoff = 1.640609780e-08 pvoff = -3.279393560e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.968798717e+00 lnfactor = -1.643739784e-05 wnfactor = -3.312238968e-07 pnfactor = 6.620791413e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.128410307e-02 lu0 = -2.074325610e-07 wu0 = -5.732509211e-09 pu0 = 1.145863814e-13
+ ua = 1.368212397e-09 lua = -4.335209226e-14 wua = -1.330909162e-15 pua = 2.660337022e-20
+ ub = 1.679787904e-19 lub = 2.487685152e-23 wub = 8.973976729e-25 pub = -1.793796542e-29
+ uc = -1.117224743e-10 luc = 1.211222431e-16 wuc = 4.137206980e-18 puc = -8.269809248e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.421845430e+05 lvsat = -1.239880483e+00 wvsat = -2.888185426e-02 pvsat = 5.773156301e-7
+ a0 = 2.078607149e+00 la0 = -1.228530240e-05 wa0 = -2.651577759e-07 pa0 = 5.300204312e-12
+ ags = 1.426154198e-01 lags = -5.861820045e-07 wags = -1.749214772e-08 pags = 3.496482668e-13
+ a1 = 0.0
+ a2 = 1.522317962e+00 la2 = -1.104021193e-05 wa2 = -2.571713939e-07 pa2 = 5.140565560e-12
+ b0 = -3.733154313e-07 lb0 = 5.406698123e-12 wb0 = 8.814776441e-14 pb0 = -1.761974204e-18
+ b1 = -6.753716816e-07 lb1 = 1.354624695e-11 wb1 = 3.974997031e-13 pb1 = -7.945569890e-18
+ keta = 7.873486781e-02 lketa = -1.106855868e-06 wketa = -2.610002932e-08 pketa = 5.217100931e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.880260953e-01 lpclm = 8.056036225e-06 wpclm = 1.869131312e-07 ppclm = -3.736182281e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 9.024796093e-03 lpdiblc2 = -1.548665147e-07 wpdiblc2 = -4.168393459e-09 ppdiblc2 = 8.332147496e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 4.384806970e+08 lpscbe1 = 7.226362351e+03 wpscbe1 = 2.117136573e+02 ppscbe1 = -4.231916773e-3
+ pscbe2 = 3.320298000e-09 lpscbe2 = 1.347315202e-13 wpscbe2 = 3.247657028e-15 ppscbe2 = -6.491699414e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.248929186e-10 lalpha0 = 6.494242313e-15 walpha0 = 1.512772905e-16 palpha0 = -3.023862094e-21
+ alpha1 = -3.248929186e-10 lalpha1 = 6.494242313e-15 walpha1 = 1.512772905e-16 palpha1 = -3.023862094e-21
+ beta0 = 1.177210880e+02 lbeta0 = -1.753445424e-03 wbeta0 = -4.084486844e-05 pbeta0 = 8.164427654e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.359282047e-09 lagidl = -2.916425399e-14 wagidl = -3.228354500e-16 pagidl = 6.453115841e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.432067107e-01 lkt1 = 4.096853045e-06 wkt1 = 1.164460877e-07 pkt1 = -2.327625709e-12
+ kt2 = -7.467703956e-02 lkt2 = 3.224412527e-07 wkt2 = 5.553115523e-09 pkt2 = -1.110005043e-13
+ at = -5.657680575e+04 lat = 2.549916296e+00 wat = 7.830376234e-02 pat = -1.565203726e-6
+ ute = 5.912473887e-01 lute = -1.347704362e-05 wute = -1.854629326e-08 pute = 3.707194450e-13
+ ua1 = 6.134683819e-09 lua1 = -8.084466128e-14 wua1 = -1.385827039e-15 pua1 = 2.770111652e-20
+ ub1 = -5.657513470e-18 lub1 = 8.852297894e-23 wub1 = 1.765490015e-24 pub1 = -3.529015039e-29
+ uc1 = -1.323423940e-10 luc1 = 2.049926460e-15 wuc1 = 2.235391544e-17 puc1 = -4.468295096e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.182 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.001190484e+00 lvth0 = -9.789475491e-08 wvth0 = -3.958482110e-08 pvth0 = 7.782740030e-14
+ k1 = 5.348733406e-01 lk1 = 3.271326537e-08 wk1 = -4.364197099e-08 pk1 = -5.115496977e-14
+ k2 = 2.688621804e-02 lk2 = -1.410272908e-07 wk2 = -6.736157027e-09 pk2 = 8.417784970e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.374102039e-01 lvoff = 2.053264710e-07 wvoff = -1.807863175e-08 pvoff = -5.244533475e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -3.361767208e-01 lnfactor = 9.965621291e-06 wnfactor = 8.596922930e-07 pnfactor = -2.893283208e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = -1.858285159e-02 lu0 = 1.110593572e-07 wu0 = 1.604451965e-08 pu0 = -5.938747115e-14
+ ua = -7.304475204e-09 lua = 2.593288153e-14 wua = 3.780973236e-15 pua = -1.423479372e-20
+ ub = 5.184541336e-18 lub = -1.519981451e-23 wub = -2.418352441e-24 pub = 8.551131192e-30
+ uc = -8.496157175e-11 luc = -9.266712812e-17 wuc = -1.291118286e-17 puc = 5.349927763e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.958154602e+04 lvsat = 6.915573731e-01 wvsat = 9.545760975e-02 pvsat = -4.160161837e-7
+ a0 = -2.386114571e-01 la0 = 6.226655804e-06 wa0 = 8.247078741e-07 pa0 = -3.406590684e-12
+ ags = -5.369205286e-03 lags = 5.960479275e-07 wags = 2.971107168e-08 pags = -2.745211655e-14
+ a1 = 0.0
+ a2 = -5.174269096e-01 la2 = 5.255044677e-06 wa2 = 7.715141817e-07 pa2 = -3.077469774e-12
+ b0 = 5.128059880e-07 lb0 = -1.672410700e-12 wb0 = -2.652318605e-13 pb0 = 1.061129681e-18
+ b1 = 2.022462712e-06 lb1 = -8.006401306e-12 wb1 = -1.184928410e-12 pb1 = 4.696242589e-18
+ keta = -9.938390274e-02 lketa = 3.161118346e-07 wketa = 6.261515623e-08 pketa = -1.870239913e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.897111865e-01 lpclm = 1.126504620e-05 wpclm = 2.246038229e-07 ppclm = -4.037288317e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.054616505e-02 lpdiblc2 = 8.137204970e-08 wpdiblc2 = 1.216857279e-08 ppdiblc2 = -4.719242458e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1.884557909e+09 lpscbe1 = -4.326160507e+03 wpscbe1 = -6.351409718e+02 ppscbe1 = 2.533494768e-3
+ pscbe2 = 3.302779523e-08 lpscbe2 = -1.025978132e-13 wpscbe2 = -1.078530388e-14 ppscbe2 = 4.719050623e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 9.746787557e-10 lalpha0 = -3.887866848e-15 walpha0 = -4.538318716e-16 palpha0 = 1.810276338e-21
+ alpha1 = 9.746787557e-10 lalpha1 = -3.887866848e-15 walpha1 = -4.538318716e-16 palpha1 = 1.810276338e-21
+ beta0 = -2.331632640e+02 lbeta0 = 1.049724049e-03 wbeta0 = 1.225346053e-04 pbeta0 = -4.887746111e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.273818749e-09 lagidl = -2.848149881e-14 wagidl = -1.511223337e-15 pagidl = 1.594699218e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.832074918e-01 lkt1 = -3.304149585e-06 wkt1 = -4.082542109e-07 pkt1 = 1.864136765e-12
+ kt2 = -1.015288132e-02 lkt2 = -1.930338593e-07 wkt2 = -1.665934657e-08 pkt2 = 6.645196775e-14
+ at = 3.076922906e+05 lat = -3.601821589e-01 wat = -1.669313473e-01 pat = 3.939476842e-7
+ ute = -1.773777213e+00 lute = 5.416830465e-06 wute = -8.032099971e-08 pute = 8.642295441e-13
+ ua1 = -1.004325146e-08 lua1 = 4.839876052e-14 wua1 = 4.157481117e-15 pua1 = -1.658365170e-20
+ ub1 = 1.195721866e-17 lub1 = -5.219882614e-23 wub1 = -5.296470045e-24 pub1 = 2.112693047e-29
+ uc1 = 2.167821799e-09 luc1 = -1.632578625e-14 wuc1 = -9.470643324e-16 puc1 = 7.297726848e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.183 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.058219043e+00 lvth0 = 1.295847556e-07 wvth0 = -3.084764775e-09 pvth0 = -6.776657936e-14
+ k1 = 4.420413699e-01 lk1 = 4.030079283e-07 wk1 = -3.259001331e-08 pk1 = -9.523979222e-14
+ k2 = 1.244243493e-02 lk2 = -8.341291769e-08 wk2 = 1.471276377e-08 pk2 = -1.379106991e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.583304515e-01 ldsub = -1.190001388e-06 wdsub = 2.259675247e-14 pdsub = -9.013550883e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.516497707e-01 lvoff = 2.621262519e-07 wvoff = 2.029611000e-09 pvoff = -1.326545010e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 9.485268245e-01 lnfactor = 4.841105860e-06 wnfactor = 7.364477754e-07 pnfactor = -2.401676849e-12
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391132325e-01 letab = 2.756836997e-7
+ u0 = 1.327885685e-02 lu0 = -1.603285579e-08 wu0 = -1.160052684e-09 pu0 = 9.239331286e-15
+ ua = -3.069262731e-09 lua = 9.039169554e-15 wua = 1.566218255e-15 pua = -5.400424015e-21
+ ub = 6.031517940e-18 lub = -1.857829408e-23 wub = -3.002336697e-24 pub = 1.088056847e-29
+ uc = -8.830803216e-11 luc = -7.931853261e-17 wuc = -2.638083478e-17 puc = 1.072279681e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.787700283e+05 lvsat = -4.187508712e-01 wvsat = -5.581668455e-02 pvsat = 1.873973106e-7
+ a0 = 1.823564999e+00 la0 = -1.999097994e-06 wa0 = -2.488887635e-07 pa0 = 8.758467362e-13
+ ags = -6.119319565e-01 lags = 3.015547889e-06 wags = 3.346854552e-07 pags = -1.243955286e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.500816326e-07 lb0 = 9.717618431e-13 wb0 = 1.320779002e-13 pb0 = -5.236873045e-19
+ b1 = 9.645726915e-08 lb1 = -3.238159745e-13 wb1 = -5.283617142e-14 pb1 = 1.804738219e-19
+ keta = 2.476080193e-04 lketa = -8.130530974e-08 wketa = 1.305224933e-08 pketa = 1.067600116e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.759158628e+00 lpclm = -2.890934136e-06 wpclm = -1.260104079e-06 ppclm = 1.885018491e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -7.745269496e-04 lpdiblc2 = 2.505555624e-09 wpdiblc2 = 6.988029947e-10 ppdiblc2 = -1.441003946e-15
+ pdiblcb = -1.195605023e+00 lpdiblcb = 3.871617257e-06 wpdiblcb = 4.519350518e-07 ppdiblcb = -1.802710170e-12
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 4.818903939e-09 lpscbe2 = 9.923786967e-15 wpscbe2 = 2.283964872e-15 ppscbe2 = -4.941107795e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.944350000e-11 lalpha0 = 3.966671938e-16
+ alpha1 = -9.944350000e-11 lalpha1 = 3.966671938e-16
+ beta0 = 5.062987286e+01 lbeta0 = -8.228988095e-05 wbeta0 = 2.147046717e-06 pbeta0 = -8.564290239e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.170570912e-09 lagidl = 1.213203773e-15 wagidl = 2.403884430e-15 pagidl = 3.301362624e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.578050196e-01 lkt1 = 1.646087992e-06 wkt1 = 3.057690869e-07 pkt1 = -9.840093464e-13
+ kt2 = -5.655244364e-02 lkt2 = -7.952037149e-09 wkt2 = -3.852746317e-09 pkt2 = 1.536810420e-14
+ at = 2.778422636e+05 lat = -2.411142819e-01 wat = -6.807471536e-02 pat = -3.785691357e-10
+ ute = -3.615564910e+00 lute = 1.276348216e-05 wute = 2.062825386e-06 pute = -7.684502778e-12
+ ua1 = -3.949854351e-10 lua1 = 9.913081626e-15 wua1 = 1.913990138e-15 pua1 = -7.634657842e-21
+ ub1 = -1.544915052e-18 lub1 = 1.659429959e-24 wub1 = -2.029866285e-25 pub1 = 8.096872730e-31
+ uc1 = -3.810527422e-09 luc1 = 7.521071603e-15 wuc1 = 1.722458408e-15 puc1 = -3.350652326e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.184 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.039402605e+00 lvth0 = 9.216130506e-08 wvth0 = -2.437274475e-08 pvth0 = -2.542755462e-14
+ k1 = 6.750746429e-01 lk1 = -6.046495744e-08 wk1 = -9.872576197e-08 pk1 = 3.629561422e-14
+ k2 = -2.822260898e-02 lk2 = -2.535431808e-09 wk2 = 1.345277469e-08 pk2 = 1.126847487e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.099377798e+00 ldsub = -5.647153224e-06 wdsub = -1.662802093e-06 pdsub = 3.307097154e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.667254791e-01 lvoff = 9.322287599e-08 wvoff = -3.305072519e-08 pvoff = -6.288427276e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.762524345e+00 lnfactor = 1.233300612e-06 wnfactor = -2.090695125e-07 pnfactor = -5.211658803e-13
+ eta0 = -1.519541026e+00 leta0 = 3.023163996e-06 weta0 = 6.066980445e-07 peta0 = -1.206643540e-12
+ etab = -3.242478655e+00 letab = 6.447874088e-06 wetab = 1.899006599e-06 petab = -3.776877255e-12
+ u0 = 7.322833509e-03 lu0 = -4.187099650e-09 wu0 = 3.193370718e-09 pu0 = 5.809380853e-16
+ ua = 1.219224695e-09 lua = 5.099255679e-16 wua = -8.772250411e-16 pua = -5.407329460e-22
+ ub = -2.684319370e-18 lub = -1.243626726e-24 wub = 2.060338836e-24 pub = 8.115649823e-31
+ uc = -2.517262462e-10 luc = 2.456990507e-16 wuc = 7.811128004e-17 puc = -1.005932643e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.587901898e+05 lvsat = 2.526125199e-01 wvsat = 1.023597558e-01 pvsat = -1.271950663e-7
+ a0 = -1.052230102e-01 la0 = 1.837010613e-06 wa0 = 6.676304502e-07 pa0 = -9.469908324e-13
+ ags = 2.157354643e+00 lags = -2.492203149e-06 wags = -1.115236789e-06 pags = 1.639751569e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 4.352185734e-07 lb0 = -1.923241775e-13 wb0 = -1.833554166e-13 pb0 = 1.036685563e-19
+ b1 = 1.727920353e-08 lb1 = -1.663410951e-13 wb1 = -1.748716152e-14 pb1 = 1.101692366e-19
+ keta = -1.290819922e-01 lketa = 1.759144522e-07 wketa = 6.550315553e-08 pketa = -9.364203266e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.107973809e+00 lpclm = 3.930578153e-07 wpclm = -1.130567811e-07 ppclm = -3.963094679e-13
+ pdiblc1 = 4.121363472e-01 lpdiblc1 = -4.402631691e-08 wpdiblc1 = -9.685305112e-09 ppdiblc1 = 1.926281278e-14
+ pdiblc2 = 5.399081098e-04 lpdiblc2 = -1.086848325e-10 wpdiblc2 = -5.117563388e-11 ppdiblc2 = 5.060604908e-17
+ pdiblcb = 1.716210045e+00 lpdiblcb = -1.919604377e-06 wpdiblcb = -9.038701037e-07 ppdiblcb = 8.938100294e-13
+ drout = 8.015169287e-01 ldrout = -4.803457740e-07 wdrout = -2.435715807e-07 pdrout = 4.844322098e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.015329920e-08 lpscbe2 = -6.856317339e-16 wpscbe2 = -2.307566904e-16 ppscbe2 = 6.034647795e-23
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.134202365e-11 lalpha0 = 1.763291894e-16 walpha0 = 5.192006143e-17 palpha0 = -1.032622526e-22
+ alpha1 = -6.673993786e-10 lalpha1 = 1.526257602e-15 walpha1 = 4.494059589e-16 palpha1 = -8.938100294e-22
+ beta0 = 1.119916002e+01 lbeta0 = -3.867319100e-06 wbeta0 = -3.820958616e-06 pbeta0 = 3.305296529e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.840433132e-09 lagidl = 1.050095265e-14 wagidl = 5.426532653e-15 pagidl = -5.681518111e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.763963195e-01 lkt1 = -8.085780255e-07 wkt1 = -4.119049211e-07 pkt1 = 4.433509579e-13
+ kt2 = -8.325143714e-02 lkt2 = 4.514879005e-08 wkt2 = 1.405519212e-08 pkt2 = -2.024845732e-14
+ at = 2.142530865e+05 lat = -1.146436752e-01 wat = -1.088087953e-01 pat = 8.063622035e-8
+ ute = 6.757041188e+00 lute = -7.866282934e-06 wute = -3.668456273e-06 pute = 3.714271374e-12
+ ua1 = 8.872030529e-09 lua1 = -8.517808414e-15 wua1 = -3.429118983e-15 pua1 = 2.992091596e-21
+ ub1 = -1.093224513e-18 lub1 = 7.610761966e-25 wub1 = -2.764821611e-25 pub1 = 9.558603327e-31
+ uc1 = 3.050590158e-11 luc1 = -1.182443435e-16 wuc1 = -1.523980640e-17 puc1 = 1.054035220e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.185 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.393630562e-01 lvth0 = -6.764803059e-09 wvth0 = -6.522320028e-08 pvth0 = 1.496823534e-14
+ k1 = 1.036233135e+00 lk1 = -4.176037558e-07 wk1 = -2.674904405e-07 pk1 = 2.031819418e-13
+ k2 = -2.039832981e-01 lk2 = 1.712690408e-07 wk2 = 9.838001200e-08 pk2 = -8.285514968e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -8.949702736e+00 ldsub = 6.267821044e-06 wdsub = 4.969690856e-06 pdsub = -3.251576149e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 5.508940289e-02 lvoff = -1.261232064e-07 wvoff = -1.674328432e-07 pvoff = 7.000217228e-14
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -3.452426112e+00 lnfactor = 7.379078670e-06 wnfactor = 2.252107746e-06 pnfactor = -2.954950236e-12
+ eta0 = 4.861051927e+00 leta0 = -3.286412958e-06 weta0 = -2.283895339e-06 peta0 = 1.651777539e-12
+ etab = 6.487716274e+00 letab = -3.174023772e-06 wetab = -3.800221049e-06 petab = 1.858917989e-12
+ u0 = -6.391795367e-02 lu0 = 6.626077757e-08 wu0 = 3.515284552e-08 pu0 = -3.102282776e-14
+ ua = -6.591124033e-09 lua = 8.233345115e-15 wua = 2.363224143e-15 pua = -3.745115931e-21
+ ub = -8.487567513e-18 lub = 4.495031265e-24 wub = 5.066304269e-24 pub = -2.160944055e-30
+ uc = 1.576238271e-10 luc = -1.590949563e-16 wuc = -1.151140133e-16 puc = 9.048143153e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.116220372e+05 lvsat = -1.479001907e-02 wvsat = -3.938743769e-02 pvsat = 1.297448089e-8
+ a0 = 1.344493545e+00 la0 = 4.034294024e-07 wa0 = 3.073766263e-08 pa0 = -3.171866615e-13
+ ags = -1.939894728e+00 lags = 1.559443836e-06 wags = 1.073854730e-06 pags = -5.249753618e-13
+ a1 = 0.0
+ a2 = 2.913840811e+00 la2 = -2.090313763e-06 wa2 = -1.061644519e-06 pa2 = 1.049828416e-12
+ b0 = 4.761008263e-07 lb0 = -2.327514109e-13 wb0 = -1.552922291e-13 pb0 = 7.591771203e-20
+ b1 = -2.985084183e-07 lb1 = 1.459318104e-13 wb1 = 1.857534144e-13 pb1 = -9.080927169e-20
+ keta = 1.935815657e-01 lketa = -1.431578603e-07 wketa = -8.964129099e-08 pketa = 5.977565617e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.061344774e+00 lpclm = 4.391678689e-07 wpclm = -1.417790393e-07 ppclm = -3.679068884e-13
+ pdiblc1 = 4.431003231e-01 lpdiblc1 = -7.464566375e-08 wpdiblc1 = 1.456474821e-07 ppdiblc1 = -1.343411205e-13
+ pdiblc2 = -2.882175809e-03 lpdiblc2 = 3.275311292e-09 wpdiblc2 = 1.725747505e-09 ppdiblc2 = -1.706539935e-15
+ pdiblcb = 2.488695745e-01 lpdiblcb = -4.685954062e-07 wpdiblcb = -2.775084480e-07 ppdiblcb = 2.744197790e-13
+ drout = 1.975396214e+00 ldrout = -1.641159782e-06 wdrout = -5.971208369e-07 pdrout = 8.340464627e-13
+ pscbe1 = 3.957407796e+09 lpscbe1 = -3.122265847e+03 wpscbe1 = -1.470158533e+03 ppscbe1 = 1.453795668e-3
+ pscbe2 = -3.195998947e-07 lpscbe2 = 3.253974091e-13 wpscbe2 = 1.530238043e-13 ppscbe2 = -1.514884912e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.773159527e-10 lalpha0 = -8.668444980e-17 walpha0 = -1.038401229e-16 palpha0 = 5.076432086e-23
+ alpha1 = 1.634798757e-09 lalpha1 = -7.503170684e-16 walpha1 = -8.988119177e-16 palpha1 = 4.394021822e-22
+ beta0 = 5.113065223e+00 lbeta0 = 2.151037458e-06 wbeta0 = -3.330506028e-07 pbeta0 = -1.437910686e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.951882136e-09 lagidl = -1.160114153e-15 wagidl = -8.223340539e-16 pagidl = 4.977987103e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.732833718e-01 lkt1 = 1.305317309e-07 wkt1 = 1.164958543e-07 pkt1 = -7.916871696e-14
+ kt2 = -1.613356663e-02 lkt2 = -2.122205856e-08 wkt2 = -1.269939897e-08 pkt2 = 6.208355176e-15
+ at = 1.162303488e+05 lat = -1.771193063e-02 wat = -5.392306603e-02 pat = 2.636136929e-8
+ ute = -1.870039733e+00 lute = 6.647785763e-07 wute = 1.776831840e-08 pute = 6.907446245e-14
+ ua1 = -2.421503566e-09 lua1 = 2.650028647e-15 wua1 = -3.411093850e-17 pua1 = -3.651300094e-22
+ ub1 = 4.668020406e-19 lub1 = -7.815872610e-25 wub1 = 1.212877246e-24 pub1 = -5.169225039e-31
+ uc1 = -1.103061339e-10 luc1 = 2.100045407e-17 wuc1 = 1.806666692e-16 puc1 = -8.832251459e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.186 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.026208119e+00 lvth0 = 3.569114285e-08 wvth0 = 1.890568325e-08 pvth0 = -2.615985195e-14
+ k1 = 8.188028463e-01 lk1 = -3.113086104e-07 wk1 = -3.047637114e-07 pk1 = 2.214037258e-13
+ k2 = -1.553872427e-01 lk2 = 1.475118872e-07 wk2 = 1.268195278e-07 pk2 = -9.675837577e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.366663739e+00 ldsub = -1.219891035e-06 wdsub = -3.022304140e-06 pdsub = 6.554704447e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -6.648274296e-01 lvoff = 2.258225355e-07 wvoff = 2.480315105e-07 pvoff = -1.331058863e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.191062040e+01 lnfactor = -5.020153877e-06 wnfactor = -8.721049739e-06 pnfactor = 2.409497264e-12
+ eta0 = -4.108147213e+00 leta0 = 1.098359425e-06 weta0 = 2.140998501e-06 peta0 = -5.114203123e-13
+ etab = -9.184020961e-03 letab = 2.115875312e-09 wetab = 4.273372071e-09 petab = -9.851980944e-16
+ u0 = 1.225082940e-01 lu0 = -2.487742213e-08 wu0 = -4.952951183e-08 pu0 = 1.037583628e-14
+ ua = 1.904840340e-08 lua = -4.301050663e-15 wua = -9.180321284e-15 pua = 1.898177122e-21
+ ub = 5.498519906e-19 lub = 7.690799229e-26 wub = 7.966673929e-25 pub = -7.364667538e-32
+ uc = -3.225775581e-10 luc = 7.566109490e-17 wuc = 1.341133172e-16 puc = -3.135833352e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.210888892e+05 lvsat = -1.941807899e-02 wvsat = -4.623513880e-02 pvsat = 1.632211653e-8
+ a0 = 5.696410685e+00 la0 = -1.724092330e-06 wa0 = -2.404335403e-06 pa0 = 8.732475082e-13
+ ags = 5.810000578e-02 lags = 5.826841502e-07 wags = 5.549748591e-07 pags = -2.713105594e-13
+ a1 = 0.0
+ a2 = -4.697481834e+00 la2 = 1.630633538e-06 wa2 = 2.869137901e-06 pa2 = -8.718131861e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.510404719e-01 lketa = 2.531751523e-08 wketa = 5.632197244e-08 pketa = -1.158140442e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.925681103e+00 lpclm = -9.611202324e-07 wpclm = -2.160216954e-06 ppclm = 6.188468548e-13
+ pdiblc1 = -6.227259153e-01 lpdiblc1 = 4.464048094e-07 wpdiblc1 = 2.182871636e-07 ppdiblc1 = -1.698524816e-13
+ pdiblc2 = -7.707258018e-03 lpdiblc2 = 5.634149232e-09 wpdiblc2 = 6.348467793e-10 ppdiblc2 = -1.173231298e-15
+ pdiblcb = -8.788827743e-01 lpdiblcb = 8.272888460e-08 wpdiblcb = 4.181909030e-07 ppdiblcb = -6.568676277e-14
+ drout = -1.466578777e+00 ldrout = 4.151853117e-08 wdrout = 1.149336726e-06 pdrout = -1.974424604e-14
+ pscbe1 = -5.514807670e+09 lpscbe1 = 1.508416128e+03 wpscbe1 = 2.940327369e+03 ppscbe1 = -7.023585744e-4
+ pscbe2 = 6.699202243e-07 lpscbe2 = -1.583492914e-13 wpscbe2 = -3.077454202e-13 ppscbe2 = 7.376775954e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.073916704e+01 lbeta0 = -5.993949375e-07 wbeta0 = -1.606972851e-06 pbeta0 = 4.789913008e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.197358382e-08 lagidl = -5.570553456e-15 wagidl = -5.966871468e-15 pagidl = 3.012808716e-21
+ bgidl = -1.179124819e+08 lbgidl = 5.465138750e+02 wbgidl = 5.205246456e+02 pbgidl = -2.544688835e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.624250724e-01 lkt1 = -2.143756591e-08 wkt1 = -4.929672926e-08 pkt1 = 1.882303386e-15
+ kt2 = -2.712052184e-02 lkt2 = -1.585086577e-08 wkt2 = -2.275412971e-08 pkt2 = 1.112381139e-14
+ at = 2.293166184e+05 lat = -7.299641525e-02 wat = -8.066565581e-02 pat = 3.943501915e-8
+ ute = 1.318134179e+00 lute = -8.938240039e-07 wute = -5.781723559e-07 pute = 3.604119799e-13
+ ua1 = 5.576685961e-09 lua1 = -1.260046268e-15 wua1 = -1.523518861e-15 pua1 = 3.629968418e-22
+ ub1 = -1.221665322e-18 lub1 = 4.385377850e-26 wub1 = -1.820449962e-25 pub1 = 1.650131326e-31
+ uc1 = 1.084614330e-10 luc1 = -8.594844639e-17 wuc1 = -8.587146652e-17 puc1 = 4.197998384e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.187 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 7.352342750e-02 lvth0 = -2.270017317e-07 wvth0 = -5.330968799e-07 pvth0 = 1.056970003e-13
+ k1 = -6.298412839e+00 lk1 = 1.388780700e-06 wk1 = 3.329223700e-06 pk1 = -6.466468472e-13
+ k2 = 2.782500184e+00 lk2 = -5.542612823e-07 wk2 = -1.358652162e-06 pk2 = 2.580762468e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.387487042e+00 ldsub = -9.859950972e-07 wdsub = -2.200227547e-06 pdsub = 4.591010091e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 2.055226571e+00 lvoff = -4.239167637e-07 wvoff = -1.135527989e-06 pvoff = 1.973849713e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -7.492669133e+00 lnfactor = 2.003409893e-06 wnfactor = 5.271201214e-06 pnfactor = -9.328317212e-13
+ eta0 = 4.900000037e-01 leta0 = -2.509388253e-16 weta0 = -1.704107522e-15 peta0 = 1.168426467e-22
+ etab = 8.855911077e-03 letab = -2.193323254e-09 wetab = -4.126417165e-09 petab = 1.021259560e-15
+ u0 = 6.609382791e-02 lu0 = -1.140169861e-08 wu0 = -2.831732711e-08 pu0 = 5.308881712e-15
+ ua = 1.238063328e-08 lua = -2.708320415e-15 wua = -6.513081556e-15 pua = 1.261053568e-21
+ ub = -3.346776898e-18 lub = 1.007695735e-24 wub = 2.452625144e-24 pub = -4.692053034e-31
+ uc = 1.394789572e-10 luc = -3.471034490e-17 wuc = -6.482432146e-17 puc = 1.616190021e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.114884930e+05 lvsat = -6.489883236e-02 wvsat = -1.044099100e-01 pvsat = 3.021832412e-8
+ a0 = -4.600347823e+00 la0 = 7.354943751e-07 wa0 = 2.685085077e-06 pa0 = -3.424623619e-13
+ ags = 5.506785593e+00 lags = -7.188433760e-07 wags = -1.982053021e-06 pags = 3.347092904e-13
+ a1 = 0.0
+ a2 = 2.686163724e+00 la2 = -1.330978760e-07 wa2 = -1.040044856e-06 pa2 = 6.197329922e-14
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700592797e-01 lketa = 5.374753786e-08 wketa = 1.126062763e-07 pketa = -2.502603607e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.549166851e-02 lpclm = -4.620288215e-08 wpclm = 3.404477442e-07 ppclm = 2.151307839e-14
+ pdiblc1 = 1.829534444e+00 lpdiblc1 = -1.393666226e-07 wpdiblc1 = -7.644425520e-07 ppdiblc1 = 6.489216557e-14
+ pdiblc2 = 1.022867181e-01 lpdiblc2 = -2.064011184e-08 wpdiblc2 = -4.450988237e-08 ppdiblc2 = 9.610490155e-15
+ pdiblcb = 9.486856462e+00 lpdiblcb = -2.393335247e-06 wpdiblcb = -4.522054030e-06 ppdiblcb = 1.114389544e-12
+ drout = -6.841647336e+00 ldrout = 1.325461158e-06 wdrout = 3.650360836e-06 pdrout = -6.171638752e-13
+ pscbe1 = 7.996773148e+08 lpscbe1 = 7.509940378e-02 wpscbe1 = 1.356055240e-01 ppscbe1 = -3.496793459e-8
+ pscbe2 = 5.045485777e-08 lpscbe2 = -1.037759935e-14 wpscbe2 = -1.915446704e-14 ppscbe2 = 4.832038563e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.477571885e+01 lbeta0 = -1.563606069e-06 wbeta0 = -2.649624018e-06 pbeta0 = 7.280493850e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.351758246e-08 lagidl = 2.907221434e-15 wagidl = 1.231284124e-14 pagidl = -1.353666259e-21
+ bgidl = 4.992544064e+09 lbgidl = -6.742208802e+02 wbgidl = -1.859016352e+03 pbgidl = 3.139320747e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.989131219e-01 lkt1 = -1.794114204e-07 wkt1 = -3.911379023e-07 pkt1 = 8.353790439e-14
+ kt2 = -1.173440897e-01 lkt2 = 5.700837883e-09 wkt2 = 3.492681360e-08 pkt2 = -2.654435537e-15
+ at = 5.077620567e+05 lat = -1.395086771e-01 wat = -1.875157839e-01 pat = 6.495830924e-8
+ ute = -6.560091088e+00 lute = 9.880476656e-07 wute = 2.856619414e-06 pute = -4.600567301e-13
+ ua1 = -3.452041285e-10 lua1 = 1.545156182e-16 wua1 = 2.973155380e-16 pua1 = -7.194587116e-23
+ ub1 = -1.690910674e-18 lub1 = 1.559424157e-25 wub1 = 8.127360648e-25 pub1 = -7.261021949e-32
+ uc1 = -1.058809044e-09 luc1 = 1.928774524e-16 wuc1 = 4.658427252e-16 puc1 = -8.980798513e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.188 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -2.561522121e+00 lvth0 = 2.399221122e-07 wvth0 = 6.999056940e-07 pvth0 = -1.128407605e-13
+ k1 = 5.014142124e+00 lk1 = -5.740765128e-07 wk1 = -2.229347261e-06 pk1 = 3.214273464e-13
+ k2 = -1.747039533e+00 lk2 = 2.318472505e-07 wk2 = 8.997322661e-07 pk2 = -1.357093495e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.070246770e-01 ldsub = 1.035850396e-08 wdsub = 9.683496291e-07 pdsub = -8.362512053e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -3.281552362e+00 lvoff = 5.253549948e-07 wvoff = 1.377137027e-06 pvoff = -2.497734971e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 5.105877086e+01 lnfactor = -8.677864679e-06 wnfactor = -2.283980411e-05 pnfactor = 4.198253458e-12
+ eta0 = 7.760982113e+00 leta0 = -1.351457445e-06 weta0 = -3.385529233e-06 peta0 = 6.292683184e-13
+ etab = 3.959197557e-01 letab = -7.435768005e-08 wetab = -1.828549683e-07 petab = 3.434434469e-14
+ u0 = 3.808276950e-02 lu0 = -7.343082539e-09 wu0 = -1.625333523e-08 pu0 = 3.600988171e-15
+ ua = 1.156351902e-09 lua = -8.947075586e-16 wua = -1.390286124e-15 pua = 4.358287769e-22
+ ub = 6.970520919e-18 lub = -8.085365335e-25 wub = -2.625559720e-24 pub = 4.274424163e-31
+ uc = -7.672994775e-10 luc = 1.303383017e-16 wuc = 4.043708594e-16 puc = -6.942040324e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.189746534e+05 lvsat = 1.201000421e-01 wvsat = 4.436449237e-01 pvsat = -6.860657469e-8
+ a0 = -6.935358078e+00 la0 = 1.243544328e-06 wa0 = 4.162627355e-06 pa0 = -6.515685413e-13
+ ags = 1.250000270e+00 lags = -4.235737183e-14 wags = -1.255811632e-13 pags = 1.972252406e-20
+ a1 = 0.0
+ a2 = 7.693463499e-01 la2 = 2.097821188e-07 wa2 = -5.869303230e-07 pa2 = -1.600829949e-14
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.001720002e+00 lketa = 1.951520354e-07 wketa = 4.267164202e-07 pketa = -8.592903841e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.285013399e+00 lpclm = 7.633503896e-07 wpclm = 2.869001892e-06 ppclm = -4.463035776e-13
+ pdiblc1 = 5.165122340e+00 lpdiblc1 = -7.733822648e-07 wpdiblc1 = -2.258240345e-06 ppdiblc1 = 3.490770007e-13
+ pdiblc2 = -1.049004960e-01 lpdiblc2 = 1.579195305e-08 wpdiblc2 = 5.919108705e-08 ppdiblc2 = -8.696929121e-15
+ pdiblcb = -3.668849702e+01 lpdiblcb = 5.948342671e-06 wpdiblcb = 1.765861111e-05 ppdiblcb = -2.896146032e-12
+ drout = 1.045574033e+00 ldrout = -7.103624891e-09 wdrout = -2.668906125e-08 pdrout = 4.160024129e-15
+ pscbe1 = 1.259780903e+09 lpscbe1 = -8.543679443e+01 wpscbe1 = -2.141737918e+02 ppscbe1 = 3.979519955e-5
+ pscbe2 = -1.104974066e-07 lpscbe2 = 1.849389388e-14 wpscbe2 = 5.541536989e-14 ppscbe2 = -8.541819795e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -7.893512919e-02 lbeta0 = 1.040021567e-06 wbeta0 = 5.968381082e-06 pbeta0 = -8.004871074e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.441165268e-08 lagidl = -9.426117981e-15 wagidl = -2.225190933e-14 pagidl = 4.934611494e-21
+ bgidl = 1.000001312e+09 lbgidl = -2.042606182e-04 wbgidl = -6.108383255e-04 pbgidl = 9.510823774e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.227239905e-01 lkt1 = 1.100607382e-08 wkt1 = 8.520428022e-08 pkt1 = 3.409873068e-15
+ kt2 = 7.944095580e-01 lkt2 = -1.631929141e-07 wkt2 = -3.740163109e-07 pkt2 = 7.308860324e-14
+ at = -2.609334921e+06 lat = 4.258219176e-01 wat = 1.428116186e+00 pat = -2.287999070e-7
+ ute = -3.545751960e+00 lute = 5.272383744e-07 wute = 8.196532909e-07 pute = -1.277593586e-13
+ ua1 = 1.536643681e-09 lua1 = -1.797084777e-16 wua1 = -1.910596230e-15 pua1 = 3.311959592e-22
+ ub1 = -1.057100144e-18 lub1 = 5.383464358e-26 wub1 = 2.172518994e-24 pub1 = -3.326626819e-31
+ uc1 = -4.085983784e-11 luc1 = 2.308804341e-17 wuc1 = 5.102270534e-17 puc1 = -2.174628191e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.189 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.0909503
+ k1 = 0.43165561
+ k2 = 0.019248026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.26995672
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.1464712
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0109067
+ ua = -8.0059916e-10
+ ub = 1.41251395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.0283e-7
+ b1 = 2.3178e-9
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.190 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.099880192e+00 lvth0 = 1.784984565e-7
+ k1 = 4.317673477e-01 lk1 = -2.233509594e-9
+ k2 = 2.048102620e-02 lk2 = -2.464628068e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.116597486e-06 lcit = 1.287534022e-10 wcit = -1.482307658e-27 pcit = -2.032879073e-32
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.734999503e-01 lvoff = 7.082516944e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.257440798e+00 lnfactor = -2.218156878e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.972594573e-03 lu0 = 3.866058195e-8
+ ua = -1.490134421e-09 lua = 1.378303069e-14
+ ub = 2.095288224e-18 lub = -1.364788619e-23
+ uc = -1.028371403e-10 luc = -5.648554281e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.509137115e+00 la0 = -9.022399339e-07 wa0 = -8.881784197e-22
+ ags = 1.050481491e-01 lags = 1.647452859e-7
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.840035766e-07 lb0 = 1.622568070e-12
+ b1 = 1.783244563e-07 lb1 = -3.518174171e-12 wb1 = -3.474158573e-29 pb1 = 9.264422861e-35
+ keta = 2.268075241e-02 lketa = 1.360255782e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.340066551e-02 lpclm = 3.196888926e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 7.248400546e-05 lpdiblc2 = 2.408008786e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.931706757e+08 lpscbe1 = -1.862376525e+3
+ pscbe2 = 1.029517683e-08 lpscbe2 = -4.688425941e-15 wpscbe2 = 6.617444900e-30
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.665939700e-09 lagidl = -1.530512396e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.931195419e-01 lkt1 = -9.021068602e-7
+ kt2 = -6.275080858e-02 lkt2 = 8.404937201e-8
+ at = 1.115934318e+05 lat = -8.116167193e-1
+ ute = 5.514161667e-01 lute = -1.268086250e-05 wute = -5.551115123e-23
+ ua1 = 3.158391808e-09 lua1 = -2.135194718e-14 pua1 = 1.323488980e-35
+ ub1 = -1.865832633e-18 lub1 = 1.273156360e-23 pub1 = -6.162975822e-45
+ uc1 = -8.433367566e-11 luc1 = 1.090286431e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.191 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.086205412e+00 lvth0 = 6.925241662e-8
+ k1 = 4.411450137e-01 lk1 = -7.715046481e-8
+ k2 = 1.241921041e-02 lk2 = 3.975851759e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.762370458e-01 lvoff = 9.269146934e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.510154194e+00 lnfactor = 3.751818661e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.587539919e-02 lu0 = -1.648502680e-8
+ ua = 8.157880917e-10 lua = -4.638684493e-15
+ ub = -9.269181748e-21 lub = 3.165149325e-24
+ uc = -1.126904653e-10 luc = 2.223138962e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.054294065e+05 lvsat = -2.019059592e-1
+ a0 = 1.532584651e+00 la0 = -1.089559245e-6
+ ags = 5.844021883e-02 lags = 5.370899819e-7
+ a1 = 0.0
+ a2 = 1.139526975e+00 la2 = -1.354328965e-6
+ b0 = -5.682315436e-08 lb0 = 6.065402102e-13 pb0 = -1.058791184e-34
+ b1 = -5.223663765e-07 lb1 = 2.079553802e-12
+ keta = 3.509246699e-02 lketa = -8.555301647e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.073374523e-01 lpclm = 2.594304016e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 5.587850927e-03 lpdiblc2 = -1.998146148e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 5.204879729e+08 lpscbe1 = 1.114937140e+3
+ pscbe2 = 9.864577265e-09 lpscbe2 = -1.248422033e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.821751706e-11 lagidl = 5.767295655e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.935857243e-01 lkt1 = 6.993914107e-7
+ kt2 = -4.593157427e-02 lkt2 = -5.031730436e-8
+ at = -5.082029532e+04 lat = 4.858854327e-01 wat = 7.275957614e-18 pat = 1.164153218e-22
+ ute = -1.946279800e+00 lute = 7.272905874e-6
+ ua1 = -1.114375423e-09 lua1 = 1.278263477e-14 pua1 = 1.654361225e-36
+ ub1 = 5.821761488e-19 lub1 = -6.825260318e-24 pub1 = -1.540743956e-45
+ uc1 = 1.338450270e-10 luc1 = -6.527148612e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.192 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.064844084e+00 lvth0 = -1.595514454e-8
+ k1 = 3.720489440e-01 lk1 = 1.984647748e-7
+ k2 = 4.404052043e-02 lk2 = -8.637477729e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.583305000e-01 ldsub = -1.190001582e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.472908466e-01 lvoff = -2.277115626e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.530169821e+00 lnfactor = -3.168910745e-7
+ eta0 = 1.590575825e-01 leta0 = -3.153504191e-7
+ etab = -1.391132325e-01 letab = 2.756836997e-7
+ u0 = 1.078745248e-02 lu0 = 3.810131197e-9
+ ua = 2.944491542e-10 lua = -2.559131245e-15
+ ub = -4.164950337e-19 lub = 4.789520309e-24
+ uc = -1.449652236e-10 luc = 1.509712047e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.889449718e+04 lvsat = -1.628425534e-2
+ a0 = 1.289035351e+00 la0 = -1.180727503e-7
+ ags = 1.068602294e-01 lags = 3.439488544e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.335774303e-07 lb0 = -1.529429699e-13
+ b1 = -1.701711870e-08 lb1 = 6.378130810e-14 wb1 = -8.271806126e-31 pb1 = 1.654361225e-36
+ keta = 2.827946504e-02 lketa = -5.837683738e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.287739745e-02 lpclm = 1.157453809e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 7.262676750e-04 lpdiblc2 = -5.892378908e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.724094998e-09 lpscbe2 = -6.880565344e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.944350000e-11 lalpha0 = 3.966671938e-16
+ alpha1 = -9.944350000e-11 lalpha1 = 3.966671938e-16
+ beta0 = 5.524100961e+01 lbeta0 = -1.006831060e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.921671662e-10 lagidl = 1.922225818e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.011155013e-01 lkt1 = -4.672342876e-7
+ kt2 = -6.482685146e-02 lkt2 = 2.505349996e-8
+ at = 1.316405906e+05 lat = -2.419273215e-1
+ ute = 8.146926502e-01 lute = -3.740254304e-06 wute = 2.220446049e-22 pute = -6.661338148e-28
+ ua1 = 3.715623896e-09 lua1 = -6.483604617e-15
+ ub1 = -1.980862298e-18 lub1 = 3.398366850e-24
+ uc1 = -1.112640540e-10 luc1 = 3.249933986e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.193 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.091747092e+00 lvth0 = 3.755143993e-8
+ k1 = 4.630447947e-01 lk1 = 1.748585722e-8
+ k2 = 6.694422700e-04 lk2 = -1.153410749e-10 wk2 = 4.336808690e-25
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.717638000e-01 ldsub = 1.455383069e-06 pdsub = -2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -2.377073596e-01 lvoff = -4.183146586e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 2.313513103e+00 lnfactor = 1.140109728e-7
+ eta0 = -2.165569650e-01 leta0 = 4.316980860e-07 weta0 = 3.035766083e-24 peta0 = 3.209238431e-29
+ etab = 8.359510565e-01 letab = -1.663592413e-06 wetab = 2.190088388e-22 petab = 1.899522206e-28
+ u0 = 1.418112353e-02 lu0 = -2.939439348e-9
+ ua = -6.647606861e-10 lua = -6.513875702e-16
+ ub = 1.740597915e-18 lub = 4.993428553e-25
+ uc = -8.396939611e-11 luc = 2.965843340e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.104425915e+04 lvsat = -2.055985244e-2
+ a0 = 1.328623436e+00 la0 = -1.968083056e-7
+ ags = -2.378002026e-01 lags = 1.029433648e-06 pags = 2.220446049e-28
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 4.143259121e-08 lb0 = 3.032113618e-14
+ b1 = -2.027735849e-08 lb1 = 7.026550122e-14
+ keta = 1.159683213e-02 lketa = -2.519724925e-08 wketa = 2.602085214e-24 pketa = -8.673617380e-31
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.651657345e-01 lpclm = -4.580820963e-07 wpclm = -4.440892099e-22
+ pdiblc1 = 3.913355579e-01 lpdiblc1 = -2.656251107e-9
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 2.784068077e-01 ldrout = 5.600522523e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.657711168e-09 lpscbe2 = -5.560277248e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.228489143e-10 lalpha0 = -4.544352013e-17
+ alpha1 = 2.977740000e-10 lalpha1 = -3.933467754e-16
+ beta0 = 2.993021526e+00 lbeta0 = 3.231350053e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.813940273e-09 lagidl = -1.701044061e-15 wagidl = 1.654361225e-30
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.082373987e-01 lkt1 = 1.435912404e-7
+ kt2 = -5.306559515e-02 lkt2 = 1.661890126e-9
+ at = -1.943173781e+04 lat = 5.853590038e-02 pat = -7.275957614e-24
+ ute = -1.121573381e+00 lute = 1.107271173e-7
+ ua1 = 1.507432243e-09 lua1 = -2.091798484e-15 pua1 = -4.135903063e-37
+ ub1 = -1.687015530e-18 lub1 = 2.813943829e-24 wub1 = 1.925929944e-40 pub1 = -5.777789833e-46
+ uc1 = -2.224094860e-12 luc1 = 1.081270951e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.194 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.079440630e+00 lvth0 = 2.538194975e-8
+ k1 = 4.617533202e-01 lk1 = 1.876295759e-8
+ k2 = 7.303995037e-03 lk2 = -6.676051270e-09 wk2 = 4.336808690e-25 pk2 = 6.505213035e-31
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.723527600e+00 ldsub = -7.154747378e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -3.045002282e-01 lvoff = 2.421799805e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 1.384346518e+00 lnfactor = 1.032835934e-6
+ eta0 = -4.398980000e-02 leta0 = 2.610515935e-7
+ etab = -1.673884872e+00 letab = 8.183090420e-7
+ u0 = 1.157857682e-02 lu0 = -3.658589740e-10
+ ua = -1.515710622e-09 lua = 1.900912925e-16
+ ub = 2.393156055e-18 lub = -1.459523120e-25
+ uc = -8.960249234e-11 luc = 3.522883326e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.703102198e+04 lvsat = 1.307481740e-2
+ a0 = 1.410507743e+00 la0 = -2.777812396e-7
+ ags = 3.663853228e-01 lags = 4.319727072e-7
+ a1 = 0.0
+ a2 = 6.337842000e-01 la2 = 1.643658181e-7
+ b0 = 1.425851653e-07 lb0 = -6.970560976e-14
+ b1 = 1.004276595e-07 lb1 = -4.909606988e-14
+ keta = 1.062116491e-03 lketa = -1.477978500e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.568509154e-01 lpclm = -3.509728211e-7
+ pdiblc1 = 7.559023000e-01 lpdiblc1 = -3.631653654e-7
+ pdiblc2 = 8.241514375e-04 lpdiblc2 = -3.897645320e-10
+ pdiblcb = -3.471255631e-01 lpdiblcb = 1.207663056e-7
+ drout = 6.929807845e-01 ldrout = 1.500924839e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.043950024e-09 lpscbe2 = 5.090225685e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.430217145e-11 lalpha0 = 2.234029744e-17
+ alpha1 = -2.955480000e-10 lalpha1 = 1.933715508e-16
+ beta0 = 4.397784152e+00 lbeta0 = 1.842222435e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.185784198e-09 lagidl = -9.100936318e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.230893210e-01 lkt1 = -3.949613924e-8
+ kt2 = -4.340761934e-02 lkt2 = -7.888592413e-9
+ at = 4.216756200e+02 lat = 3.890345544e-2
+ ute = -1.831879340e+00 lute = 8.131273709e-7
+ ua1 = -2.494762429e-09 lua1 = 1.865851762e-15 wua1 = 8.271806126e-31 pua1 = -4.135903063e-37
+ ub1 = 3.071655861e-18 lub1 = -1.891763550e-24 pub1 = 7.703719778e-46
+ uc1 = 2.777053201e-10 luc1 = -1.686867054e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.195 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -9.856050479e-01 lvth0 = -2.049145151e-8
+ k1 = 1.642725377e-01 lk1 = 1.641923878e-7
+ k2 = 1.169785987e-01 lk2 = -6.029267476e-08 wk2 = 2.775557562e-23 pk2 = 6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.242326091e-01 ldsub = 1.878397956e-07 pdsub = 5.551115123e-29
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -1.321388743e-01 lvoff = -6.004429701e-8
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.180728471e+00 lnfactor = 1.546386882e-7
+ eta0 = 0.49
+ etab = -6.25e-6
+ u0 = 1.613550270e-02 lu0 = -2.593603331e-9
+ ua = -6.678498755e-10 lua = -2.244023905e-16
+ ub = 2.260826543e-18 lub = -8.126038331e-26 wub = -1.540743956e-39
+ uc = -3.454710167e-11 luc = 8.313904430e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.179130700e+04 lvsat = 1.563635687e-2
+ a0 = 5.327040663e-01 la0 = 1.513506437e-7
+ ags = 1.25
+ a1 = 0.0
+ a2 = 1.464464770e+00 la2 = -2.417289920e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.007975172e-02 lketa = 4.445401076e-10
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.137409036e-01 lpclm = 3.679554014e-07 wpclm = 2.775557562e-23 ppclm = 5.551115123e-29
+ pdiblc1 = -1.539182482e-01 lpdiblc1 = 8.161860606e-08 wpdiblc1 = -2.775557562e-23 ppdiblc1 = -1.040834086e-29
+ pdiblc2 = -6.343819909e-03 lpdiblc2 = 3.114441620e-09 wpdiblc2 = 7.318364664e-25 ppdiblc2 = -5.624298770e-31
+ pdiblcb = 1.925112622e-02 lpdiblcb = -5.834426652e-8
+ drout = 1.001811303e+00 ldrout = -8.854919108e-10
+ pscbe1 = 8.000300498e+08 lpscbe1 = -1.469046821e-2
+ pscbe2 = 8.986204433e-09 lpscbe2 = 7.913234404e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.287927943e+00 lbeta0 = 4.293178398e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.412562592e-10 lagidl = 8.999499052e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.682979248e-01 lkt1 = -1.739500910e-8
+ kt2 = -7.598876628e-02 lkt2 = 8.039352891e-9
+ at = 5.607382532e+04 lat = 1.169678902e-2
+ ute = 7.641373640e-02 lute = -1.197798653e-07 pute = -2.775557562e-29
+ ua1 = 2.304678064e-09 lua1 = -4.804507120e-16
+ ub1 = -1.612636960e-18 lub1 = 3.982466821e-25
+ uc1 = -7.596169672e-11 luc1 = 4.210489046e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.196 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = 5.565e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = -1.07139
+ k1 = 0.85164386
+ k2 = -0.1354293
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.66213569
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = -0.38350697
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = 3.8281044
+ eta0 = 0.49
+ etab = -6.25e-6
+ u0 = 0.0052777
+ ua = -1.607283e-9
+ ub = 1.9206399e-18
+ uc = 2.58041e-13
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 87251.0
+ a0 = 1.166315
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.45249595
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.028218739
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.82665932
+ pdiblc1 = 0.18776805
+ pdiblc2 = 0.0066944085
+ pdiblcb = -0.225
+ drout = 0.9981043
+ pscbe1 = 799968550.0
+ pscbe2 = 9.3174823e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.0852145
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.9262738e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.4765e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.54112
+ kt2 = -0.042333
+ at = 105041.0
+ ute = -0.42503
+ ua1 = 2.9333e-10
+ ub1 = 5.4574e-20
+ uc1 = -5.8335e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.197 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre)
+ toxe = 4.01004e-09
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -2.2811e-8
+ lint = -2.935e-9
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre)
+ vth0 = 1.830266384e+00 lvth0 = -5.393308720e-07 wvth0 = -1.345007653e-06 pvth0 = 2.499965725e-13
+ k1 = -1.747554175e+00 lk1 = 4.831129388e-07 wk1 = 9.190472936e-07 pk1 = -1.708233205e-13
+ k2 = 1.560235661e-01 lk2 = -5.417234423e-08 wk2 = 1.362421986e-08 pk2 = -2.532333746e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.670698446e+00 ldsub = -1.116811559e-06 wdsub = -2.373756167e-06 pdsub = 4.412100587e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre)
+ voff = 4.695605026e+00 lvoff = -9.440545467e-07 wvoff = -2.337202950e-06 pvoff = 4.344159124e-13
*(mismatch parameter sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre)
+ nfactor = -3.699298928e+01 lnfactor = 7.587416682e-06 wnfactor = 1.815903255e-05 pnfactor = -3.375219380e-12
+ eta0 = 8.182383703e+00 leta0 = -1.429783359e-06 weta0 = -3.581743085e-06 peta0 = 6.657385871e-13
+ etab = 4.457253357e-01 letab = -8.284812984e-08 wetab = -2.060455421e-07 petab = 3.829768491e-14
+ u0 = -9.592712154e-02 lu0 = 1.881094018e-08 wu0 = 4.614461826e-08 pu0 = -8.576900196e-15
+ ua = -1.721190682e-08 lua = 2.900431429e-15 wua = 7.162379237e-15 pua = -1.331271429e-21
+ ub = -6.442381324e-18 lub = 1.554434755e-24 wub = 3.619782649e-24 pub = -6.728090009e-31
+ uc = -3.828960618e-10 luc = 7.121685309e-17 wuc = 2.253841722e-16 puc = -4.189215609e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.439234038e+06 lvsat = -2.512930872e-01 wvsat = -5.612645236e-01 pvsat = 1.043222370e-7
+ a0 = 1.797062686e+00 la0 = -1.172370724e-07 wa0 = 9.662013410e-08 pa0 = -1.795878433e-14
+ ags = 1.249999985e+00 lags = 2.731505688e-15 wags = 6.842682865e-15 pags = -1.271849293e-21
+ a1 = 0.0
+ a2 = -8.632484378e+00 la2 = 1.688625294e-06 wa2 = 3.790768904e-06 pa2 = -7.045902162e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.555859553e+00 lketa = 2.839425980e-07 wketa = 6.847359863e-07 pketa = -1.272718778e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.943877222e+00 lpclm = -2.076572915e-07 wpclm = -3.130661704e-08 ppclm = 5.818960909e-15
+ pdiblc1 = 9.440897930e-02 lpdiblc1 = 1.735265047e-08 wpdiblc1 = 1.027953514e-07 ppdiblc1 = -1.910657197e-14
+ pdiblc2 = 6.230151542e-02 lpdiblc2 = -1.033569296e-08 wpdiblc2 = -1.866184791e-08 ppdiblc2 = 3.468677671e-15
+ pdiblcb = -9.647124730e+00 lpdiblcb = 1.751290324e-06 wpdiblcb = 5.067553259e-06 ppdiblcb = -9.419061243e-13
+ drout = 9.882548598e-01 ldrout = 1.830715458e-09 wdrout = 6.956739185e-15 pdrout = -1.293049223e-21
+ pscbe1 = 1.285433399e+09 lpscbe1 = -9.023335140e+01 wpscbe1 = -2.261181578e+02 ppscbe1 = 4.202858199e-5
+ pscbe2 = 1.576995002e-08 lpscbe2 = -1.199320176e-15 wpscbe2 = -3.377489220e-15 ppscbe2 = 6.277739214e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.257026038e+01 lbeta0 = -2.506465477e-06 wbeta0 = -4.577582627e-06 pbeta0 = 8.508352829e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.487813614e-07 lagidl = 2.819789816e-14 wagidl = 6.770300827e-14 pagidl = -1.258395815e-20
+ bgidl = 1.000000010e+09 lbgidl = -1.901000977e-06 wbgidl = -4.762187958e-06 pbgidl = 8.851480484e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 6.265e-9
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 5.46384e-11
+ cgdo = 5.46384e-11
+ cgbo = 0.0
+ cgdl = 6.920864e-12
+ cgsl = 6.920864e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000672644022
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.60458928e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.299366688e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 6.243816758e-01 lkt1 = -2.166317965e-07 wkt1 = -5.885999544e-07 pkt1 = 1.094030735e-13
+ kt2 = 1.111362601e+00 lkt2 = -2.144374014e-07 wkt2 = -5.215966208e-07 pkt2 = 9.694916391e-14
+ at = -1.175221209e+04 lat = 2.170835433e-02 wat = 2.186245303e-01 pat = -4.063574145e-8
+ ute = -1.785411394e+00 lute = 2.528540896e-07 wute = -4.483453608e-15 pute = 8.333396195e-22
+ ua1 = -3.768870207e-11 lua1 = 6.152644615e-17 wua1 = -1.177552437e-15 pua1 = 2.188716715e-22
+ ub1 = 4.060735096e-18 lub1 = -7.446251629e-25 wub1 = -2.104576860e-25 pub1 = 3.911777010e-32
+ uc1 = -9.759609062e-10 luc1 = 1.705591272e-16 wuc1 = 4.864263350e-16 puc1 = -9.041206288e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
