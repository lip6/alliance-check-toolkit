../rtl/cla16.vhdl