* Pad_15800W12000H
.subckt Pad_15800W12000H pad

.ends Pad_15800W12000H
