* BulkConn_4000WNoUp
* BulkConn_4000WNoUp
.subckt BulkConn_4000WNoUp vdd vss iovdd iovss

.ends BulkConn_4000WNoUp
