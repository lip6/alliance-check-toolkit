* Spice description of oa2ao222_x4
* Spice driver version -1162834149
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:34

* INTERF i0 i1 i2 i3 i4 q vdd vss 


.subckt oa2ao222_x4 10 11 7 5 6 4 3 13 
* NET 3 = vdd
* NET 4 = q
* NET 5 = i3
* NET 6 = i4
* NET 7 = i2
* NET 10 = i0
* NET 11 = i1
* NET 13 = vss
Mtr_00014 3 9 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 4 9 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 2 5 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 1 7 9 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 9 6 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 2 11 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 3 10 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 4 9 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 13 9 4 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 8 5 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00004 12 10 13 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00003 9 11 12 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00002 8 6 9 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00001 13 7 8 13 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
C12 2 13 9.75335e-16
C11 3 13 4.04764e-15
C10 4 13 2.20321e-15
C9 5 13 1.50967e-15
C8 6 13 1.376e-15
C7 7 13 1.52801e-15
C6 8 13 4.67807e-16
C5 9 13 2.96334e-15
C4 10 13 1.69828e-15
C3 11 13 1.38512e-15
C1 13 13 4.23938e-15
.ends oa2ao222_x4

