* PNP_05v5_W0u68L0u68
.subckt PNP_05v5_W0u68L0u68 collector base emitter
Xpnp collector base emitter sky130_fd_pr__pnp_05v5_W0p68L0p68
.ends PNP_05v5_W0u68L0u68
