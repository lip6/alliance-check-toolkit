* Spice description of xr2_x4
* Spice driver version -15180005
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:45

* INTERF i0 i1 q vdd vss 


.subckt xr2_x4 9 4 3 2 10 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i1
* NET 9 = i0
* NET 10 = vss
Mtr_00016 2 8 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 3 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 8 4 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 1 11 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 2 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 5 4 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00010 2 9 11 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 1 9 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 5 4 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00007 10 8 3 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 3 8 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 6 11 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 8 5 7 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 10 4 6 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 10 9 11 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 7 9 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C11 1 10 1.19992e-15
C10 2 10 4.91083e-15
C9 3 10 2.15173e-15
C8 4 10 2.44863e-15
C7 5 10 2.05671e-15
C4 8 10 3.2943e-15
C3 9 10 2.54824e-15
C2 10 10 3.30621e-15
C1 11 10 1.66447e-15
.ends xr2_x4

