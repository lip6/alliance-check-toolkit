* deprecated C4M.Sky130 global lib file
* Use the C4M.Sky130_all_lib.spice instead
.lib tt
.include "C4M.Sky130_logic_tt_model.spice"
.include "C4M.Sky130_io_tt_model.spice"
.include "C4M.Sky130_diode_tt_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl tt
.lib ff
.include "C4M.Sky130_logic_ff_model.spice"
.include "C4M.Sky130_io_ff_model.spice"
.include "C4M.Sky130_diode_ff_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl ff
.lib ss
.include "C4M.Sky130_logic_ss_model.spice"
.include "C4M.Sky130_io_ss_model.spice"
.include "C4M.Sky130_diode_ss_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl ss
.lib fs
.include "C4M.Sky130_logic_fs_model.spice"
.include "C4M.Sky130_io_fs_model.spice"
.include "C4M.Sky130_diode_fs_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl fs
.lib sf
.include "C4M.Sky130_logic_sf_model.spice"
.include "C4M.Sky130_io_sf_model.spice"
.include "C4M.Sky130_diode_sf_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl sf
