-- no model for and21nor_x1
