* SP6TCell
.subckt SP6TCell vdd vss wl bl bl_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 bit_n bit vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 bit_n bit vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl wl bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg2 bl_n wl bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
.ends SP6TCell
