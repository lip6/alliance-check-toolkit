* dffnr_x1
.subckt dffnr_x1 vdd vss i clk q nrst
Mclk_nmos _clk_n clk vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_pmos _clk_n clk vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos0 vss _clk_n _clk_buf vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos0 vdd _clk_n _clk_buf vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi_nmos _u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi_pmos _u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mu_nmos vss _u _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mu_pmos vdd _u _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos1 _net0 _clk_n _dff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_buf_pmos0 _net1 _clk_buf _dff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_buf_nmos0 _dff_m _clk_buf _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos1 _dff_m _clk_n _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
My_nmos _net2 _y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
My_pmos _net3 _y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mdff_m_nmos vss _dff_m _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mdff_m_pmos vdd _dff_m _y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_nmos0 _net6 nrst _y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnrst_pmos0 _y nrst vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_pmos1 vdd nrst _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mclk_buf_nmos1 _y _clk_buf _dff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_nmos2 _dff_s _clk_n _net7 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_n_pmos2 _y _clk_n _dff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mnrst_nmos1 _net7 nrst _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mclk_buf_pmos1 _dff_s _clk_buf _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mq_nmos _net4 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mq_pmos _net5 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mdff_s_nmos vss _dff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.925um
Mdff_s_pmos vdd _dff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.485um
.ends dffnr_x1
