* Filler1000
.subckt Filler1000 vss vdd iovss iovdd

.ends Filler1000
