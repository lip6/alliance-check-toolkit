* Filler4000
* Filler4000
.subckt Filler4000 vss vdd iovss iovdd

.ends Filler4000
