../rtl/alu16.vhdl