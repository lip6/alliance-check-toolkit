-- no model for fill_w4
