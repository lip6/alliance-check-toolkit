* Spice description of on12_x4
* Spice driver version 433499931
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:38

* INTERF i0 i1 q vdd vss 


.subckt on12_x4 6 4 3 2 7 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i1
* NET 6 = i0
* NET 7 = vss
Mtr_00010 2 4 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00009 3 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 2 5 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 8 5 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00006 2 6 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 7 6 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 7 5 3 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 3 5 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 7 4 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 5 8 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C7 2 7 2.86631e-15
C6 3 7 2.15173e-15
C5 4 7 2.28354e-15
C4 5 7 2.18376e-15
C3 6 7 2.33846e-15
C2 7 7 2.51079e-15
C1 8 7 1.67373e-15
.ends on12_x4

