* Spice description of a2_x2
* Spice driver version 28367784
* Date ( dd/mm/yyyy hh:mm:ss ): 17/07/2024 at  8:36:49

* INTERF i0 i1 q vdd vss 


.subckt a2_x2 1 2 4 3 7 
* NET 1 = i0
* NET 2 = i1
* NET 3 = vdd
* NET 4 = q
* NET 7 = vss
Mtr_00006 4 5 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.8U AS=0.784P AD=0.784P PS=6.16U PD=6.16U 
Mtr_00005 5 1 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.4U AS=0.392P AD=0.392P PS=3.36U PD=3.36U 
Mtr_00004 3 2 5 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.4U AS=0.392P AD=0.392P PS=3.36U PD=3.36U 
Mtr_00003 7 5 4 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.4U AS=0.392P AD=0.392P PS=3.36U PD=3.36U 
Mtr_00002 6 2 5 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.4U AS=0.392P AD=0.392P PS=3.36U PD=3.36U 
Mtr_00001 7 1 6 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.4U AS=0.392P AD=0.392P PS=3.36U PD=3.36U 
C7 1 7 8.8444e-16
C6 2 7 1.18445e-15
C5 3 7 1.60117e-15
C4 4 7 1.36257e-15
C3 5 7 1.96274e-15
C1 7 7 1.56724e-15
.ends a2_x2

