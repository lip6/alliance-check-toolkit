* Filler200
.subckt Filler200 vss vdd iovss iovdd

.ends Filler200
