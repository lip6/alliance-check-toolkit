* Spice description of rowend_x0
* Spice driver version -262557925
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:30:04

* INTERF vdd vss 


.subckt rowend_x0 1 2 
* NET 1 = vdd
* NET 2 = vss
C2 1 2 3.8726e-16
C1 2 2 3.8726e-16
.ends rowend_x0

