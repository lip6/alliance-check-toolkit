* xor2_x0
.subckt xor2_x0 vdd vss i0 i1 q
Mi0_nmos0 i0_n i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos0 i0_n i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_nmos1 vss i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_pmos1 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos0 _net0 i1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_n_pmos _net1 i1_n q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi0_n_nmos q i0_n _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi0_n_pmos q i0_n _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_n_nmos _net2 i1_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos0 _net1 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mi1_nmos1 vss i1 i1_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mi1_pmos1 vdd i1 i1_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends xor2_x0
