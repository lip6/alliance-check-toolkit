* Spice description of arlet6502_cts_r
* Spice driver version -874538072
* Date ( dd/mm/yyyy hh:mm:ss ):  7/06/2024 at  1:08:56

* INTERF a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] a[9] a[10] a[11] a[12] 
* INTERF a[13] a[14] a[15] clk di[0] di[1] di[2] di[3] di[4] di[5] di[6] 
* INTERF di[7] do[0] do[1] do[2] do[3] do[4] do[5] do[6] do[7] irq nmi rdy 
* INTERF reset vdd vss we 


.subckt arlet6502_cts_r 2182 1530 1978 1490 1525 1474 3300 3063 2390 8156 8136 8109 8089 8066 8038 8015 4022 8055 7970 7803 6987 6804 6485 5880 4712 2502 1742 1753 1306 7406 6466 5833 4929 4230 1699 4079 3792 8144 8185 1368 
* NET 65 = subckt_1739_sff1_x4.sff_s
* NET 67 = subckt_1739_sff1_x4.y
* NET 69 = subckt_1739_sff1_x4.sff_m
* NET 70 = subckt_1739_sff1_x4.u
* NET 71 = subckt_1739_sff1_x4.ckr
* NET 72 = subckt_1739_sff1_x4.nckr
* NET 73 = subckt_1622_sff1_x4.sff_s
* NET 75 = subckt_1622_sff1_x4.y
* NET 76 = subckt_1622_sff1_x4.sff_m
* NET 79 = subckt_1622_sff1_x4.u
* NET 80 = subckt_1622_sff1_x4.ckr
* NET 81 = subckt_1622_sff1_x4.nckr
* NET 83 = subckt_1623_sff1_x4.sff_s
* NET 85 = subckt_1623_sff1_x4.y
* NET 87 = subckt_1623_sff1_x4.sff_m
* NET 88 = subckt_1623_sff1_x4.u
* NET 89 = subckt_1623_sff1_x4.ckr
* NET 90 = subckt_1623_sff1_x4.nckr
* NET 91 = abc_11867_auto_rtlil_cc_2608_muxgate_11616
* NET 96 = subckt_1637_sff1_x4.sff_s
* NET 99 = subckt_1637_sff1_x4.y
* NET 100 = subckt_1637_sff1_x4.sff_m
* NET 101 = subckt_1637_sff1_x4.u
* NET 103 = subckt_1637_sff1_x4.ckr
* NET 104 = subckt_1637_sff1_x4.nckr
* NET 106 = subckt_1650_sff1_x4.sff_s
* NET 107 = subckt_1650_sff1_x4.y
* NET 110 = subckt_1650_sff1_x4.sff_m
* NET 111 = subckt_1650_sff1_x4.u
* NET 112 = subckt_1650_sff1_x4.ckr
* NET 113 = subckt_1650_sff1_x4.nckr
* NET 115 = subckt_1632_sff1_x4.sff_s
* NET 116 = subckt_1632_sff1_x4.y
* NET 119 = subckt_1632_sff1_x4.sff_m
* NET 120 = subckt_1632_sff1_x4.u
* NET 121 = subckt_1632_sff1_x4.ckr
* NET 122 = subckt_1632_sff1_x4.nckr
* NET 123 = subckt_1647_sff1_x4.sff_s
* NET 125 = subckt_1647_sff1_x4.y
* NET 126 = subckt_1647_sff1_x4.sff_m
* NET 129 = subckt_1647_sff1_x4.u
* NET 130 = subckt_1647_sff1_x4.ckr
* NET 131 = subckt_1647_sff1_x4.nckr
* NET 133 = subckt_1617_sff1_x4.sff_s
* NET 134 = subckt_1617_sff1_x4.y
* NET 137 = subckt_1617_sff1_x4.sff_m
* NET 138 = subckt_1617_sff1_x4.u
* NET 139 = subckt_1617_sff1_x4.ckr
* NET 140 = subckt_1617_sff1_x4.nckr
* NET 141 = abc_11867_auto_rtlil_cc_2608_muxgate_11604
* NET 146 = subckt_1631_sff1_x4.sff_s
* NET 148 = subckt_1631_sff1_x4.y
* NET 149 = subckt_1631_sff1_x4.sff_m
* NET 152 = subckt_1631_sff1_x4.u
* NET 153 = subckt_1631_sff1_x4.ckr
* NET 154 = subckt_1631_sff1_x4.nckr
* NET 159 = abc_11867_new_n872
* NET 161 = abc_11867_new_n871
* NET 163 = abc_11867_new_n877
* NET 165 = abc_11867_new_n878
* NET 166 = abc_11867_new_n860
* NET 169 = subckt_1655_sff1_x4.sff_s
* NET 170 = subckt_1655_sff1_x4.y
* NET 173 = subckt_1655_sff1_x4.sff_m
* NET 174 = subckt_1655_sff1_x4.u
* NET 175 = subckt_1655_sff1_x4.ckr
* NET 176 = subckt_1655_sff1_x4.nckr
* NET 177 = abc_11867_auto_rtlil_cc_2608_muxgate_11670
* NET 185 = abc_11867_new_n608
* NET 187 = abc_11867_new_n1175
* NET 190 = mos6502_nmi_1
* NET 192 = subckt_1656_sff1_x4.sff_s
* NET 193 = subckt_1656_sff1_x4.y
* NET 196 = subckt_1656_sff1_x4.sff_m
* NET 197 = subckt_1656_sff1_x4.u
* NET 198 = subckt_1656_sff1_x4.ckr
* NET 199 = subckt_1656_sff1_x4.nckr
* NET 248 = subckt_1653_sff1_x4.sff_s
* NET 249 = subckt_1653_sff1_x4.y
* NET 250 = subckt_1653_sff1_x4.sff_m
* NET 253 = subckt_1653_sff1_x4.ckr
* NET 254 = subckt_1653_sff1_x4.u
* NET 255 = subckt_1653_sff1_x4.nckr
* NET 256 = abc_11867_auto_rtlil_cc_2608_muxgate_11664
* NET 261 = abc_11867_auto_rtlil_cc_2608_muxgate_11614
* NET 266 = mos6502_axys_2_6
* NET 268 = mos6502_axys_3_6
* NET 272 = abc_11867_auto_rtlil_cc_2608_muxgate_11632
* NET 273 = mos6502_axys_0_6
* NET 278 = subckt_1648_sff1_x4.sff_s
* NET 280 = subckt_1648_sff1_x4.y
* NET 282 = subckt_1648_sff1_x4.sff_m
* NET 284 = subckt_1648_sff1_x4.u
* NET 285 = subckt_1648_sff1_x4.ckr
* NET 286 = subckt_1648_sff1_x4.nckr
* NET 287 = abc_11867_auto_rtlil_cc_2608_muxgate_11654
* NET 292 = abc_11867_auto_rtlil_cc_2608_muxgate_11622
* NET 298 = subckt_1634_sff1_x4.sff_s
* NET 299 = subckt_1634_sff1_x4.y
* NET 302 = subckt_1634_sff1_x4.sff_m
* NET 303 = subckt_1634_sff1_x4.ckr
* NET 304 = subckt_1634_sff1_x4.u
* NET 305 = subckt_1634_sff1_x4.nckr
* NET 306 = abc_11867_auto_rtlil_cc_2608_muxgate_11652
* NET 312 = subckt_1649_sff1_x4.sff_s
* NET 313 = subckt_1649_sff1_x4.y
* NET 316 = subckt_1649_sff1_x4.sff_m
* NET 317 = subckt_1649_sff1_x4.ckr
* NET 318 = subckt_1649_sff1_x4.u
* NET 319 = subckt_1649_sff1_x4.nckr
* NET 320 = abc_11867_auto_rtlil_cc_2608_muxgate_11620
* NET 325 = subckt_1633_sff1_x4.sff_s
* NET 327 = subckt_1633_sff1_x4.y
* NET 329 = subckt_1633_sff1_x4.sff_m
* NET 330 = subckt_1633_sff1_x4.u
* NET 332 = subckt_1633_sff1_x4.ckr
* NET 333 = subckt_1633_sff1_x4.nckr
* NET 334 = abc_11867_new_n873
* NET 342 = abc_11867_new_n868
* NET 343 = abc_11867_new_n864
* NET 344 = abc_11867_new_n874
* NET 349 = abc_11867_new_n865
* NET 352 = abc_11867_new_n876
* NET 354 = abc_11867_new_n875
* NET 359 = abc_11867_new_n863
* NET 365 = abc_11867_new_n870
* NET 369 = abc_11867_new_n428
* NET 370 = abc_11867_new_n608_hfns_2
* NET 375 = abc_11867_new_n475
* NET 378 = abc_11867_new_n471
* NET 384 = abc_11867_new_n431_hfns_2
* NET 386 = abc_11867_new_n431
* NET 469 = subckt_1744_sff1_x4.sff_s
* NET 470 = subckt_1744_sff1_x4.y
* NET 472 = subckt_1744_sff1_x4.sff_m
* NET 474 = subckt_1744_sff1_x4.u
* NET 475 = subckt_1744_sff1_x4.ckr
* NET 476 = subckt_1744_sff1_x4.nckr
* NET 478 = subckt_1654_sff1_x4.sff_s
* NET 479 = subckt_1654_sff1_x4.y
* NET 480 = subckt_1654_sff1_x4.sff_m
* NET 483 = subckt_1654_sff1_x4.u
* NET 484 = subckt_1654_sff1_x4.ckr
* NET 485 = subckt_1654_sff1_x4.nckr
* NET 486 = subckt_1652_sff1_x4.sff_s
* NET 489 = subckt_1652_sff1_x4.y
* NET 491 = subckt_1652_sff1_x4.sff_m
* NET 492 = subckt_1652_sff1_x4.u
* NET 493 = subckt_1652_sff1_x4.ckr
* NET 494 = subckt_1652_sff1_x4.nckr
* NET 496 = abc_11867_auto_rtlil_cc_2608_muxgate_11662
* NET 497 = mos6502_axys_2_5
* NET 498 = mos6502_axys_3_5
* NET 505 = subckt_1620_sff1_x4.y
* NET 506 = subckt_1620_sff1_x4.sff_s
* NET 507 = subckt_1620_sff1_x4.sff_m
* NET 509 = subckt_1620_sff1_x4.u
* NET 510 = subckt_1620_sff1_x4.ckr
* NET 511 = subckt_1620_sff1_x4.nckr
* NET 512 = mos6502_axys_2_1
* NET 514 = mos6502_axys_0_1
* NET 517 = mos6502_axys_3_1
* NET 519 = subckt_1618_sff1_x4.sff_s
* NET 521 = subckt_1618_sff1_x4.y
* NET 523 = subckt_1618_sff1_x4.sff_m
* NET 524 = subckt_1618_sff1_x4.u
* NET 525 = subckt_1618_sff1_x4.ckr
* NET 526 = subckt_1618_sff1_x4.nckr
* NET 528 = abc_11867_auto_rtlil_cc_2608_muxgate_11606
* NET 529 = mos6502_axys_2_0
* NET 530 = mos6502_axys_3_0
* NET 532 = mos6502_axys_0_0
* NET 535 = mos6502_axys_0_2
* NET 540 = subckt_1619_sff1_x4.sff_s
* NET 541 = subckt_1619_sff1_x4.y
* NET 543 = subckt_1619_sff1_x4.sff_m
* NET 545 = subckt_1619_sff1_x4.u
* NET 546 = subckt_1619_sff1_x4.ckr
* NET 547 = subckt_1619_sff1_x4.nckr
* NET 549 = abc_11867_auto_rtlil_cc_2608_muxgate_11624
* NET 551 = abc_11867_new_n867
* NET 553 = abc_11867_new_n862
* NET 557 = abc_11867_new_n1411
* NET 558 = abc_11867_new_n857
* NET 559 = abc_11867_new_n859
* NET 562 = abc_11867_new_n476
* NET 565 = abc_11867_new_n856
* NET 568 = abc_11867_new_n475_hfns_3
* NET 574 = abc_11867_new_n490
* NET 576 = abc_11867_new_n482
* NET 579 = abc_11867_new_n430
* NET 647 = subckt_1756_sff1_x4.sff_s
* NET 648 = subckt_1756_sff1_x4.sff_m
* NET 649 = subckt_1756_sff1_x4.y
* NET 651 = subckt_1756_sff1_x4.ckr
* NET 652 = subckt_1756_sff1_x4.u
* NET 653 = subckt_1756_sff1_x4.nckr
* NET 654 = abc_11867_auto_rtlil_cc_2608_muxgate_11860
* NET 659 = abc_11867_auto_rtlil_cc_2608_muxgate_11666
* NET 664 = subckt_1624_sff1_x4.sff_s
* NET 665 = subckt_1624_sff1_x4.sff_m
* NET 666 = subckt_1624_sff1_x4.y
* NET 668 = subckt_1624_sff1_x4.ckr
* NET 669 = subckt_1624_sff1_x4.u
* NET 670 = subckt_1624_sff1_x4.nckr
* NET 671 = abc_11867_auto_rtlil_cc_2608_muxgate_11618
* NET 676 = mos6502_axys_2_7
* NET 677 = mos6502_axys_3_7
* NET 684 = subckt_1636_sff1_x4.sff_s
* NET 685 = mos6502_axys_0_5
* NET 686 = subckt_1636_sff1_x4.sff_m
* NET 688 = subckt_1636_sff1_x4.y
* NET 691 = abc_11867_auto_rtlil_cc_2608_muxgate_11630
* NET 692 = subckt_1636_sff1_x4.ckr
* NET 693 = subckt_1636_sff1_x4.u
* NET 694 = subckt_1636_sff1_x4.nckr
* NET 697 = abc_11867_auto_rtlil_cc_2608_muxgate_11658
* NET 703 = mos6502_axys_2_3
* NET 709 = mos6502_axys_0_3
* NET 710 = abc_11867_auto_rtlil_cc_2608_muxgate_11626
* NET 715 = subckt_1640_sff1_x4.sff_s
* NET 716 = subckt_1640_sff1_x4.sff_m
* NET 718 = subckt_1640_sff1_x4.y
* NET 721 = subckt_1640_sff1_x4.u
* NET 722 = subckt_1640_sff1_x4.ckr
* NET 723 = subckt_1640_sff1_x4.nckr
* NET 724 = abc_11867_auto_rtlil_cc_2608_muxgate_11656
* NET 725 = mos6502_axys_2_2
* NET 730 = subckt_1651_sff1_x4.sff_s
* NET 732 = subckt_1651_sff1_x4.sff_m
* NET 733 = subckt_1651_sff1_x4.y
* NET 736 = subckt_1651_sff1_x4.ckr
* NET 737 = subckt_1651_sff1_x4.u
* NET 738 = subckt_1651_sff1_x4.nckr
* NET 739 = mos6502_axys_3_2
* NET 740 = abc_11867_auto_rtlil_cc_2608_muxgate_11608
* NET 747 = subckt_1621_sff1_x4.sff_s
* NET 748 = subckt_1621_sff1_x4.sff_m
* NET 749 = subckt_1621_sff1_x4.y
* NET 751 = abc_11867_auto_rtlil_cc_2608_muxgate_11612
* NET 752 = subckt_1621_sff1_x4.ckr
* NET 753 = subckt_1621_sff1_x4.u
* NET 754 = subckt_1621_sff1_x4.nckr
* NET 760 = abc_11867_new_n858
* NET 762 = abc_11867_new_n1424
* NET 763 = abc_11867_new_n1410
* NET 764 = abc_11867_new_n640
* NET 774 = abc_11867_new_n380
* NET 778 = abc_11867_new_n654
* NET 782 = abc_11867_new_n471_hfns_3
* NET 786 = abc_11867_new_n482_hfns_2
* NET 791 = abc_11867_new_n473
* NET 850 = subckt_1748_sff1_x4.sff_s
* NET 851 = subckt_1748_sff1_x4.y
* NET 853 = subckt_1748_sff1_x4.sff_m
* NET 855 = subckt_1748_sff1_x4.u
* NET 856 = subckt_1748_sff1_x4.ckr
* NET 857 = subckt_1748_sff1_x4.nckr
* NET 865 = abc_11867_new_n1906
* NET 868 = subckt_1646_sff1_x4.sff_s
* NET 869 = subckt_1646_sff1_x4.y
* NET 871 = subckt_1646_sff1_x4.sff_m
* NET 873 = subckt_1646_sff1_x4.u
* NET 874 = subckt_1646_sff1_x4.ckr
* NET 875 = subckt_1646_sff1_x4.nckr
* NET 877 = subckt_1644_sff1_x4.sff_s
* NET 879 = subckt_1644_sff1_x4.y
* NET 880 = subckt_1644_sff1_x4.sff_m
* NET 882 = subckt_1644_sff1_x4.u
* NET 883 = subckt_1644_sff1_x4.ckr
* NET 884 = subckt_1644_sff1_x4.nckr
* NET 885 = abc_11867_auto_rtlil_cc_2608_muxgate_11646
* NET 890 = abc_11867_auto_rtlil_cc_2608_muxgate_11650
* NET 899 = abc_11867_auto_rtlil_cc_2608_muxgate_11610
* NET 900 = mos6502_axys_3_3
* NET 903 = abc_11867_new_n1103
* NET 907 = subckt_1642_sff1_x4.sff_s
* NET 909 = subckt_1642_sff1_x4.y
* NET 911 = subckt_1642_sff1_x4.sff_m
* NET 912 = subckt_1642_sff1_x4.u
* NET 913 = subckt_1642_sff1_x4.nckr
* NET 914 = subckt_1642_sff1_x4.ckr
* NET 915 = abc_11867_auto_rtlil_cc_2608_muxgate_11638
* NET 920 = abc_11867_auto_rtlil_cc_2608_muxgate_11660
* NET 923 = abc_11867_new_n1166
* NET 927 = subckt_1635_sff1_x4.sff_s
* NET 929 = subckt_1635_sff1_x4.y
* NET 931 = subckt_1635_sff1_x4.sff_m
* NET 932 = subckt_1635_sff1_x4.u
* NET 933 = subckt_1635_sff1_x4.ckr
* NET 934 = subckt_1635_sff1_x4.nckr
* NET 935 = abc_11867_auto_rtlil_cc_2608_muxgate_11628
* NET 939 = abc_11867_new_n1148
* NET 942 = abc_11867_new_n1421
* NET 943 = abc_11867_new_n1426
* NET 946 = abc_11867_new_n1407
* NET 947 = abc_11867_new_n1412
* NET 948 = abc_11867_new_n1409
* NET 955 = abc_11867_new_n1423
* NET 956 = abc_11867_new_n1425
* NET 957 = abc_11867_new_n663
* NET 963 = abc_11867_new_n426
* NET 965 = abc_11867_new_n490_hfns_2
* NET 969 = abc_11867_new_n430_hfns_2
* NET 1019 = subckt_1645_sff1_x4.sff_s
* NET 1020 = subckt_1645_sff1_x4.y
* NET 1022 = subckt_1645_sff1_x4.sff_m
* NET 1024 = subckt_1645_sff1_x4.u
* NET 1025 = subckt_1645_sff1_x4.nckr
* NET 1026 = subckt_1645_sff1_x4.ckr
* NET 1030 = subckt_1738_sff1_x4.sff_s
* NET 1031 = subckt_1738_sff1_x4.y
* NET 1033 = subckt_1738_sff1_x4.sff_m
* NET 1035 = subckt_1738_sff1_x4.ckr
* NET 1036 = subckt_1738_sff1_x4.u
* NET 1037 = subckt_1738_sff1_x4.nckr
* NET 1038 = abc_11867_auto_rtlil_cc_2608_muxgate_11648
* NET 1043 = mos6502_axys_1_6
* NET 1047 = abc_11867_new_n1030
* NET 1048 = mos6502_axys_1_7
* NET 1052 = abc_11867_new_n1022
* NET 1055 = subckt_1721_sff1_x4.sff_s
* NET 1056 = subckt_1721_sff1_x4.y
* NET 1058 = subckt_1721_sff1_x4.sff_m
* NET 1060 = subckt_1721_sff1_x4.u
* NET 1061 = subckt_1721_sff1_x4.ckr
* NET 1062 = subckt_1721_sff1_x4.nckr
* NET 1063 = mos6502_axys_0_7
* NET 1064 = subckt_1638_sff1_x4.sff_s
* NET 1066 = subckt_1638_sff1_x4.y
* NET 1067 = subckt_1638_sff1_x4.sff_m
* NET 1069 = abc_11867_auto_rtlil_cc_2608_muxgate_11634
* NET 1070 = subckt_1638_sff1_x4.u
* NET 1072 = subckt_1638_sff1_x4.ckr
* NET 1073 = subckt_1638_sff1_x4.nckr
* NET 1074 = abc_11867_auto_rtlil_cc_2608_muxgate_11642
* NET 1080 = subckt_1639_sff1_x4.sff_s
* NET 1081 = subckt_1639_sff1_x4.y
* NET 1083 = subckt_1639_sff1_x4.sff_m
* NET 1085 = subckt_1639_sff1_x4.ckr
* NET 1086 = subckt_1639_sff1_x4.u
* NET 1087 = subckt_1639_sff1_x4.nckr
* NET 1088 = mos6502_axys_1_1
* NET 1091 = abc_11867_auto_rtlil_cc_2608_muxgate_11636
* NET 1097 = subckt_1643_sff1_x4.sff_s
* NET 1099 = subckt_1643_sff1_x4.y
* NET 1101 = subckt_1643_sff1_x4.sff_m
* NET 1102 = subckt_1643_sff1_x4.u
* NET 1104 = subckt_1643_sff1_x4.ckr
* NET 1105 = subckt_1643_sff1_x4.nckr
* NET 1110 = abc_11867_new_n881
* NET 1111 = mos6502_axys_2_4
* NET 1113 = mos6502_axys_0_4
* NET 1114 = abc_11867_new_n882
* NET 1115 = abc_11867_new_n883
* NET 1116 = mos6502_axys_3_4
* NET 1119 = abc_11867_new_n1414
* NET 1120 = abc_11867_new_n1427
* NET 1123 = abc_11867_new_n1102
* NET 1132 = abc_11867_new_n1101
* NET 1133 = abc_11867_new_n959
* NET 1139 = abc_11867_new_n1413
* NET 1140 = abc_11867_new_n639
* NET 1145 = abc_11867_new_n1100
* NET 1148 = abc_11867_new_n766
* NET 1150 = abc_11867_new_n861
* NET 1154 = abc_11867_new_n656
* NET 1157 = abc_11867_new_n517
* NET 1167 = abc_11867_new_n606
* NET 1168 = abc_11867_new_n602
* NET 1169 = abc_11867_new_n599
* NET 1173 = abc_11867_new_n605
* NET 1184 = abc_11867_new_n426_hfns_2
* NET 1190 = abc_11867_new_n473_hfns_3
* NET 1284 = abc_11867_new_n1914
* NET 1287 = abc_11867_new_n1907
* NET 1292 = abc_11867_new_n1909
* NET 1293 = abc_11867_new_n1723
* NET 1295 = abc_11867_new_n1724
* NET 1296 = abc_11867_new_n1910
* NET 1297 = abc_11867_new_n1920
* NET 1298 = abc_11867_new_n1913
* NET 1301 = abc_11867_new_n1725
* NET 1304 = mos6502_axys_1_5
* NET 1306 = do[3]
* NET 1307 = abc_11867_auto_rtlil_cc_2608_muxgate_11790
* NET 1313 = abc_11867_new_n909
* NET 1315 = abc_11867_new_n999
* NET 1317 = mos6502_axys_1_3
* NET 1325 = abc_11867_new_n917
* NET 1327 = abc_11867_new_n914
* NET 1330 = abc_11867_auto_rtlil_cc_2608_muxgate_11644
* NET 1332 = abc_11867_new_n1157
* NET 1335 = mos6502_axys_1_4
* NET 1338 = subckt_1717_sff1_x4.sff_s
* NET 1339 = subckt_1717_sff1_x4.y
* NET 1342 = subckt_1717_sff1_x4.sff_m
* NET 1343 = subckt_1717_sff1_x4.u
* NET 1344 = subckt_1717_sff1_x4.ckr
* NET 1345 = subckt_1717_sff1_x4.nckr
* NET 1346 = abc_11867_new_n915
* NET 1348 = abc_11867_new_n916
* NET 1352 = abc_11867_new_n479
* NET 1353 = abc_11867_new_n383
* NET 1355 = abc_11867_new_n951
* NET 1356 = abc_11867_new_n1467
* NET 1357 = abc_11867_new_n1668
* NET 1358 = abc_11867_new_n1422
* NET 1359 = abc_11867_new_n1408
* NET 1361 = abc_11867_new_n1434
* NET 1362 = abc_11867_new_n855
* NET 1364 = abc_11867_new_n658
* NET 1365 = abc_11867_new_n966
* NET 1368 = we
* NET 1372 = abc_11867_new_n524
* NET 1375 = abc_11867_new_n690
* NET 1377 = abc_11867_new_n689
* NET 1381 = abc_11867_new_n641
* NET 1384 = abc_11867_new_n638
* NET 1389 = abc_11867_new_n659
* NET 1390 = abc_11867_new_n660
* NET 1446 = abc_11867_new_n1357
* NET 1451 = abc_11867_new_n1720
* NET 1455 = abc_11867_new_n1718
* NET 1466 = abc_11867_new_n1670
* NET 1467 = abc_11867_new_n1676
* NET 1473 = abc_11867_new_n1014
* NET 1474 = a[5]
* NET 1476 = abc_11867_new_n942
* NET 1477 = abc_11867_new_n943
* NET 1479 = subckt_1719_sff1_x4.sff_s
* NET 1481 = subckt_1719_sff1_x4.y
* NET 1483 = subckt_1719_sff1_x4.sff_m
* NET 1484 = subckt_1719_sff1_x4.u
* NET 1486 = subckt_1719_sff1_x4.ckr
* NET 1487 = subckt_1719_sff1_x4.nckr
* NET 1488 = abc_11867_auto_rtlil_cc_2608_muxgate_11786
* NET 1490 = a[3]
* NET 1497 = abc_11867_new_n983
* NET 1499 = mos6502_axys_1_2
* NET 1501 = subckt_1641_sff1_x4.sff_s
* NET 1502 = subckt_1641_sff1_x4.y
* NET 1504 = subckt_1641_sff1_x4.sff_m
* NET 1506 = abc_11867_auto_rtlil_cc_2608_muxgate_11640
* NET 1507 = subckt_1641_sff1_x4.ckr
* NET 1508 = subckt_1641_sff1_x4.u
* NET 1509 = subckt_1641_sff1_x4.nckr
* NET 1510 = subckt_1720_sff1_x4.sff_s
* NET 1512 = subckt_1720_sff1_x4.y
* NET 1514 = subckt_1720_sff1_x4.sff_m
* NET 1515 = subckt_1720_sff1_x4.u
* NET 1517 = subckt_1720_sff1_x4.ckr
* NET 1518 = subckt_1720_sff1_x4.nckr
* NET 1519 = abc_11867_auto_rtlil_cc_2608_muxgate_11788
* NET 1525 = a[4]
* NET 1526 = abc_11867_auto_rtlil_cc_2608_muxgate_11782
* NET 1530 = a[1]
* NET 1535 = abc_11867_new_n1420
* NET 1538 = abc_11867_new_n1417
* NET 1539 = abc_11867_new_n1415
* NET 1541 = abc_11867_new_n1418
* NET 1543 = abc_11867_new_n604
* NET 1545 = abc_11867_new_n1465
* NET 1546 = abc_11867_new_n1466
* NET 1547 = abc_11867_new_n1468
* NET 1550 = abc_11867_new_n965
* NET 1553 = abc_11867_new_n768
* NET 1558 = abc_11867_new_n1667
* NET 1559 = abc_11867_new_n598
* NET 1565 = abc_11867_new_n608_hfns_1
* NET 1570 = abc_11867_new_n509
* NET 1571 = abc_11867_new_n484
* NET 1576 = abc_11867_new_n774
* NET 1583 = abc_11867_new_n777
* NET 1587 = abc_11867_new_n613
* NET 1588 = abc_11867_new_n567
* NET 1589 = abc_11867_new_n603
* NET 1590 = abc_11867_new_n691
* NET 1593 = abc_11867_new_n580
* NET 1597 = abc_11867_new_n578
* NET 1611 = abc_11867_new_n725
* NET 1615 = abc_11867_new_n657
* NET 1616 = abc_11867_new_n652
* NET 1617 = abc_11867_new_n726
* NET 1618 = abc_11867_new_n729
* NET 1619 = abc_11867_new_n730
* NET 1621 = subckt_1630_sff1_x4.sff_s
* NET 1622 = subckt_1630_sff1_x4.y
* NET 1623 = subckt_1630_sff1_x4.sff_m
* NET 1626 = subckt_1630_sff1_x4.u
* NET 1627 = subckt_1630_sff1_x4.ckr
* NET 1628 = subckt_1630_sff1_x4.nckr
* NET 1699 = nmi
* NET 1701 = subckt_1749_sff1_x4.sff_s
* NET 1702 = subckt_1749_sff1_x4.y
* NET 1704 = subckt_1749_sff1_x4.sff_m
* NET 1706 = subckt_1749_sff1_x4.ckr
* NET 1707 = subckt_1749_sff1_x4.u
* NET 1708 = subckt_1749_sff1_x4.nckr
* NET 1710 = abc_11867_new_n1717
* NET 1711 = abc_11867_new_n1740
* NET 1719 = abc_11867_new_n1728
* NET 1727 = abc_11867_new_n1760
* NET 1729 = abc_11867_new_n1699
* NET 1732 = abc_11867_new_n1698
* NET 1738 = abc_11867_new_n927
* NET 1739 = abc_11867_new_n926
* NET 1741 = abc_11867_new_n895
* NET 1742 = do[1]
* NET 1743 = abc_11867_new_n935
* NET 1744 = abc_11867_new_n936
* NET 1746 = spare_buffer_19.q
* NET 1752 = abc_11867_new_n902
* NET 1753 = do[2]
* NET 1758 = mos6502_axys_1_0
* NET 1760 = abc_11867_new_n893
* NET 1761 = abc_11867_new_n894
* NET 1766 = subckt_1718_sff1_x4.sff_s
* NET 1767 = subckt_1718_sff1_x4.y
* NET 1768 = subckt_1718_sff1_x4.sff_m
* NET 1770 = subckt_1718_sff1_x4.u
* NET 1772 = clk_root_tr_2
* NET 1773 = subckt_1718_sff1_x4.ckr
* NET 1774 = subckt_1718_sff1_x4.nckr
* NET 1776 = abc_11867_new_n954
* NET 1778 = abc_11867_new_n953
* NET 1780 = abc_11867_new_n949
* NET 1782 = abc_11867_new_n1419
* NET 1785 = abc_11867_new_n1429
* NET 1788 = abc_11867_new_n1688
* NET 1790 = abc_11867_new_n1442
* NET 1792 = abc_11867_new_n1435
* NET 1795 = abc_11867_new_n1436
* NET 1796 = abc_11867_new_n625
* NET 1798 = abc_11867_new_n500
* NET 1799 = mos6502_state[5]
* NET 1800 = abc_11867_new_n429
* NET 1806 = abc_11867_new_n569
* NET 1807 = reset_root_tl_0
* NET 1809 = spare_buffer_14.q
* NET 1813 = abc_11867_new_n809
* NET 1816 = abc_11867_new_n830
* NET 1817 = abc_11867_new_n832
* NET 1818 = abc_11867_new_n831
* NET 1819 = abc_11867_new_n829
* NET 1821 = abc_11867_new_n775
* NET 1825 = abc_11867_new_n665
* NET 1827 = abc_11867_new_n664
* NET 1877 = subckt_1740_sff1_x4.y
* NET 1878 = subckt_1740_sff1_x4.sff_m
* NET 1887 = abc_11867_new_n583
* NET 1889 = abc_11867_new_n1437
* NET 1890 = abc_11867_new_n1441
* NET 1891 = abc_11867_new_n565
* NET 1892 = abc_11867_new_n581
* NET 1893 = abc_11867_new_n584
* NET 1897 = abc_11867_new_n644
* NET 1898 = abc_11867_new_n645
* NET 1899 = abc_11867_new_n823
* NET 1902 = abc_11867_new_n825
* NET 1904 = abc_11867_new_n525
* NET 1905 = abc_11867_new_n521
* NET 1909 = abc_11867_new_n1598
* NET 1910 = abc_11867_auto_rtlil_cc_2608_muxgate_11836
* NET 1913 = subckt_1740_sff1_x4.sff_s
* NET 1917 = subckt_1740_sff1_x4.ckr
* NET 1918 = subckt_1740_sff1_x4.u
* NET 1919 = subckt_1740_sff1_x4.nckr
* NET 1924 = abc_11867_new_n1745
* NET 1925 = abc_11867_new_n1739
* NET 1928 = abc_11867_new_n1908
* NET 1929 = abc_11867_new_n1746
* NET 1932 = abc_11867_new_n1738
* NET 1936 = abc_11867_new_n1697
* NET 1943 = abc_11867_new_n1696
* NET 1951 = clk_root_tr_1
* NET 1954 = abc_11867_new_n1912
* NET 1956 = abc_11867_new_n907
* NET 1957 = abc_11867_new_n908
* NET 1962 = abc_11867_new_n1669
* NET 1964 = abc_11867_new_n900
* NET 1965 = abc_11867_new_n901
* NET 1966 = abc_11867_new_n991
* NET 1968 = abc_11867_new_n954_hfns_2
* NET 1974 = abc_11867_auto_rtlil_cc_2608_muxgate_11784
* NET 1978 = a[2]
* NET 1985 = abc_11867_new_n1687
* NET 1986 = abc_11867_new_n530
* NET 1992 = abc_11867_new_n600
* NET 1996 = abc_11867_new_n563
* NET 1999 = abc_11867_new_n958
* NET 2003 = abc_11867_new_n1430
* NET 2005 = abc_11867_new_n1440
* NET 2006 = abc_11867_new_n850
* NET 2011 = abc_11867_new_n851
* NET 2013 = abc_11867_new_n853
* NET 2019 = spare_buffer_13.q
* NET 2022 = abc_11867_new_n776
* NET 2027 = abc_11867_new_n646
* NET 2032 = abc_11867_new_n738
* NET 2035 = abc_11867_new_n661
* NET 2036 = abc_11867_new_n666
* NET 2039 = abc_11867_new_n519
* NET 2041 = abc_11867_new_n527
* NET 2043 = abc_11867_new_n522
* NET 2126 = abc_11867_auto_rtlil_cc_2608_muxgate_11844
* NET 2127 = mos6502_alu_bi7
* NET 2132 = abc_11867_new_n1700
* NET 2133 = abc_11867_new_n1719
* NET 2135 = abc_11867_new_n1693
* NET 2136 = abc_11867_new_n1741
* NET 2138 = abc_11867_new_n1905
* NET 2141 = abc_11867_new_n1743
* NET 2143 = abc_11867_new_n1762
* NET 2144 = abc_11867_new_n1729
* NET 2152 = abc_11867_new_n1737
* NET 2154 = abc_11867_new_n1695
* NET 2155 = abc_11867_new_n1694
* NET 2156 = abc_11867_new_n1691
* NET 2159 = abc_11867_new_n1747
* NET 2166 = abc_11867_new_n1829
* NET 2167 = abc_11867_new_n1791
* NET 2168 = abc_11867_new_n1911
* NET 2170 = abc_11867_new_n1862
* NET 2172 = abc_11867_new_n885
* NET 2174 = abc_11867_new_n1816
* NET 2177 = abc_11867_new_n1817
* NET 2178 = abc_11867_new_n880
* NET 2179 = abc_11867_new_n884
* NET 2181 = abc_11867_new_n955
* NET 2182 = a[0]
* NET 2184 = subckt_1716_sff1_x4.sff_s
* NET 2185 = subckt_1716_sff1_x4.y
* NET 2188 = subckt_1716_sff1_x4.sff_m
* NET 2189 = abc_11867_auto_rtlil_cc_2608_muxgate_11780
* NET 2190 = subckt_1716_sff1_x4.u
* NET 2191 = subckt_1716_sff1_x4.ckr
* NET 2192 = subckt_1716_sff1_x4.nckr
* NET 2198 = abc_11867_new_n1039
* NET 2199 = abc_11867_new_n950
* NET 2202 = abc_11867_new_n952
* NET 2203 = abc_11867_new_n615
* NET 2205 = abc_11867_new_n1661
* NET 2206 = abc_11867_new_n1662
* NET 2207 = abc_11867_new_n1663
* NET 2210 = abc_11867_new_n579
* NET 2214 = abc_11867_new_n1689
* NET 2216 = abc_11867_new_n1439
* NET 2217 = abc_11867_new_n1438
* NET 2220 = abc_11867_new_n852
* NET 2227 = abc_11867_new_n614
* NET 2232 = abc_11867_new_n571
* NET 2233 = abc_11867_new_n566
* NET 2234 = abc_11867_new_n620
* NET 2235 = abc_11867_new_n616
* NET 2236 = abc_11867_new_n612
* NET 2238 = abc_11867_new_n834
* NET 2239 = abc_11867_new_n810
* NET 2240 = abc_11867_new_n572
* NET 2241 = abc_11867_new_n622
* NET 2242 = abc_11867_new_n817
* NET 2246 = abc_11867_new_n621
* NET 2247 = abc_11867_new_n607
* NET 2249 = abc_11867_new_n642
* NET 2251 = abc_11867_new_n650
* NET 2252 = abc_11867_new_n735
* NET 2254 = abc_11867_new_n736
* NET 2256 = abc_11867_new_n518
* NET 2258 = abc_11867_new_n516
* NET 2262 = mos6502_state[2]
* NET 2264 = subckt_1627_sff1_x4.sff_s
* NET 2265 = subckt_1627_sff1_x4.y
* NET 2267 = subckt_1627_sff1_x4.sff_m
* NET 2269 = subckt_1627_sff1_x4.u
* NET 2270 = subckt_1627_sff1_x4.ckr
* NET 2271 = subckt_1627_sff1_x4.nckr
* NET 2315 = abc_11867_new_n1026
* NET 2318 = abc_11867_new_n1722
* NET 2319 = abc_11867_auto_rtlil_cc_2608_muxgate_11846
* NET 2322 = subckt_1757_sff1_x4.sff_s
* NET 2324 = subckt_1757_sff1_x4.y
* NET 2325 = subckt_1757_sff1_x4.sff_m
* NET 2327 = subckt_1757_sff1_x4.ckr
* NET 2328 = subckt_1757_sff1_x4.u
* NET 2329 = subckt_1757_sff1_x4.nckr
* NET 2334 = abc_11867_new_n1756
* NET 2337 = abc_11867_new_n1761
* NET 2340 = abc_11867_new_n1757
* NET 2344 = abc_11867_new_n1765
* NET 2346 = abc_11867_new_n1759
* NET 2352 = abc_11867_new_n1796
* NET 2355 = abc_11867_new_n1830
* NET 2361 = abc_11867_new_n1792
* NET 2365 = abc_11867_new_n1831
* NET 2371 = abc_11867_new_n1832
* NET 2375 = abc_11867_new_n1649
* NET 2379 = abc_11867_new_n1822
* NET 2382 = abc_11867_new_n1855
* NET 2390 = a[8]
* NET 2393 = subckt_1724_sff1_x4.sff_s
* NET 2394 = subckt_1724_sff1_x4.y
* NET 2397 = subckt_1724_sff1_x4.sff_m
* NET 2398 = abc_11867_auto_rtlil_cc_2608_muxgate_11796
* NET 2399 = subckt_1724_sff1_x4.ckr
* NET 2400 = subckt_1724_sff1_x4.u
* NET 2401 = subckt_1724_sff1_x4.nckr
* NET 2402 = abc_11867_new_n1104
* NET 2407 = abc_11867_new_n961
* NET 2408 = abc_11867_new_n1046
* NET 2412 = abc_11867_new_n1041
* NET 2413 = abc_11867_new_n1044
* NET 2421 = abc_11867_new_n956
* NET 2424 = abc_11867_new_n960
* NET 2430 = abc_11867_new_n957
* NET 2437 = abc_11867_new_n1431
* NET 2439 = abc_11867_new_n1433
* NET 2441 = abc_11867_new_n1432
* NET 2448 = abc_11867_new_n724
* NET 2454 = abc_11867_new_n649
* NET 2462 = abc_11867_new_n556
* NET 2466 = abc_11867_new_n833
* NET 2467 = abc_11867_new_n835
* NET 2469 = abc_11867_new_n505
* NET 2471 = abc_11867_new_n824
* NET 2473 = abc_11867_new_n523
* NET 2477 = abc_11867_new_n800
* NET 2481 = abc_11867_new_n526
* NET 2484 = abc_11867_new_n651
* NET 2485 = abc_11867_new_n667
* NET 2490 = abc_11867_new_n485
* NET 2492 = mos6502_state[4]
* NET 2494 = subckt_1629_sff1_x4.sff_s
* NET 2495 = subckt_1629_sff1_x4.y
* NET 2496 = subckt_1629_sff1_x4.sff_m
* NET 2499 = subckt_1629_sff1_x4.ckr
* NET 2500 = subckt_1629_sff1_x4.u
* NET 2501 = subckt_1629_sff1_x4.nckr
* NET 2502 = do[0]
* NET 2589 = abc_11867_new_n1763
* NET 2591 = abc_11867_new_n1767
* NET 2594 = abc_11867_new_n1768
* NET 2595 = abc_11867_new_n1904
* NET 2596 = abc_11867_new_n1902
* NET 2599 = abc_11867_new_n1716
* NET 2601 = abc_11867_new_n1766
* NET 2602 = abc_11867_new_n1734
* NET 2605 = abc_11867_new_n1735
* NET 2608 = abc_11867_new_n1736
* NET 2610 = abc_11867_new_n1758
* NET 2612 = abc_11867_new_n1744
* NET 2614 = abc_11867_new_n1754
* NET 2616 = abc_11867_new_n1683
* NET 2619 = abc_11867_new_n1750
* NET 2621 = abc_11867_new_n1783
* NET 2630 = abc_11867_new_n1834
* NET 2631 = abc_11867_new_n1833
* NET 2635 = abc_11867_new_n1835
* NET 2636 = abc_11867_new_n1837
* NET 2638 = abc_11867_new_n1821
* NET 2642 = abc_11867_new_n1854
* NET 2648 = abc_11867_new_n1846
* NET 2652 = abc_11867_new_n1876
* NET 2659 = abc_11867_new_n1925
* NET 2661 = abc_11867_new_n1926
* NET 2663 = subckt_1750_sff1_x4.sff_s
* NET 2664 = subckt_1750_sff1_x4.y
* NET 2667 = subckt_1750_sff1_x4.sff_m
* NET 2668 = abc_11867_auto_rtlil_cc_2608_muxgate_11848
* NET 2669 = subckt_1750_sff1_x4.u
* NET 2670 = subckt_1750_sff1_x4.ckr
* NET 2671 = subckt_1750_sff1_x4.nckr
* NET 2672 = abc_11867_new_n1666
* NET 2677 = abc_11867_new_n972
* NET 2678 = abc_11867_new_n1042
* NET 2679 = abc_11867_new_n1659
* NET 2682 = abc_11867_new_n491
* NET 2687 = abc_11867_new_n382
* NET 2688 = abc_11867_new_n483
* NET 2690 = abc_11867_new_n381
* NET 2693 = abc_11867_new_n493
* NET 2695 = abc_11867_new_n767
* NET 2696 = abc_11867_new_n769
* NET 2698 = abc_11867_new_n515
* NET 2700 = abc_11867_new_n591
* NET 2702 = abc_11867_new_n590
* NET 2703 = abc_11867_new_n550
* NET 2705 = abc_11867_new_n836
* NET 2706 = abc_11867_new_n655
* NET 2707 = abc_11867_new_n506
* NET 2710 = abc_11867_new_n555
* NET 2712 = abc_11867_new_n573
* NET 2718 = abc_11867_new_n508
* NET 2719 = abc_11867_new_n653
* NET 2722 = abc_11867_new_n551
* NET 2723 = abc_11867_new_n549
* NET 2728 = subckt_1625_sff1_x4.sff_s
* NET 2729 = subckt_1625_sff1_x4.y
* NET 2732 = subckt_1625_sff1_x4.sff_m
* NET 2733 = subckt_1625_sff1_x4.u
* NET 2734 = subckt_1625_sff1_x4.ckr
* NET 2735 = subckt_1625_sff1_x4.nckr
* NET 2789 = abc_11867_new_n374
* NET 2794 = abc_11867_new_n1903
* NET 2796 = abc_11867_new_n1692
* NET 2798 = abc_11867_new_n1713
* NET 2803 = abc_11867_new_n1742
* NET 2805 = abc_11867_new_n1028
* NET 2806 = abc_11867_new_n1027
* NET 2809 = abc_11867_new_n1732
* NET 2813 = abc_11867_new_n1751
* NET 2816 = abc_11867_new_n1784
* NET 2822 = abc_11867_new_n1685
* NET 2827 = abc_11867_new_n1782
* NET 2830 = abc_11867_new_n1841
* NET 2833 = abc_11867_new_n1889
* NET 2836 = abc_11867_new_n1825
* NET 2840 = abc_11867_new_n1828
* NET 2843 = abc_11867_new_n1827
* NET 2845 = abc_11867_new_n1856
* NET 2847 = abc_11867_new_n1853
* NET 2853 = abc_11867_new_n1875
* NET 2860 = abc_11867_new_n1877
* NET 2863 = abc_11867_new_n1881
* NET 2866 = abc_11867_new_n1883
* NET 2868 = abc_11867_new_n1874
* NET 2873 = abc_11867_new_n1878
* NET 2875 = abc_11867_new_n1880
* NET 2877 = abc_11867_new_n1884
* NET 2883 = abc_11867_new_n1924
* NET 2886 = abc_11867_new_n1045
* NET 2887 = abc_11867_new_n1660
* NET 2888 = abc_11867_new_n1664
* NET 2889 = abc_11867_new_n967
* NET 2890 = abc_11867_new_n962
* NET 2894 = abc_11867_new_n499
* NET 2896 = abc_11867_new_n486
* NET 2898 = abc_11867_new_n575
* NET 2901 = abc_11867_new_n487
* NET 2904 = abc_11867_new_n770
* NET 2906 = abc_11867_new_n1428
* NET 2912 = abc_11867_new_n488
* NET 2913 = abc_11867_new_n477
* NET 2917 = abc_11867_new_n771
* NET 2918 = abc_11867_new_n701
* NET 2919 = abc_11867_new_n700
* NET 2922 = abc_11867_new_n495
* NET 2924 = abc_11867_new_n570
* NET 2925 = abc_11867_new_n806
* NET 2926 = abc_11867_new_n427
* NET 2932 = abc_11867_new_n560
* NET 2935 = abc_11867_new_n561
* NET 2937 = abc_11867_new_n763
* NET 2938 = abc_11867_new_n662
* NET 2941 = abc_11867_new_n574
* NET 2942 = abc_11867_new_n592
* NET 2943 = abc_11867_new_n562
* NET 2946 = abc_11867_new_n635
* NET 2947 = abc_11867_new_n634
* NET 2950 = abc_11867_new_n797
* NET 2951 = abc_11867_new_n798
* NET 2955 = abc_11867_new_n668
* NET 2957 = abc_11867_new_n593
* NET 2958 = abc_11867_new_n623
* NET 2961 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[5]
* NET 2962 = abc_11867_new_n837
* NET 2964 = mos6502_state[0]
* NET 2968 = mos6502_state[1]
* NET 2970 = subckt_1626_sff1_x4.sff_s
* NET 2971 = subckt_1626_sff1_x4.y
* NET 2972 = subckt_1626_sff1_x4.sff_m
* NET 2975 = subckt_1626_sff1_x4.u
* NET 2976 = subckt_1626_sff1_x4.ckr
* NET 2977 = subckt_1626_sff1_x4.nckr
* NET 3009 = abc_11867_new_n1665
* NET 3033 = abc_11867_new_n632
* NET 3063 = a[7]
* NET 3073 = abc_11867_new_n733
* NET 3077 = mos6502_pc[12]
* NET 3078 = abc_11867_new_n1024
* NET 3081 = subckt_1755_sff1_x4.sff_s
* NET 3083 = subckt_1755_sff1_x4.ckr
* NET 3084 = subckt_1755_sff1_x4.y
* NET 3085 = subckt_1755_sff1_x4.sff_m
* NET 3088 = subckt_1755_sff1_x4.u
* NET 3091 = subckt_1755_sff1_x4.nckr
* NET 3095 = abc_11867_new_n1785
* NET 3097 = abc_11867_new_n1764
* NET 3098 = abc_11867_new_n1786
* NET 3100 = abc_11867_new_n1789
* NET 3102 = abc_11867_new_n1788
* NET 3104 = abc_11867_new_n1779
* NET 3108 = abc_11867_new_n1836
* NET 3109 = abc_11867_new_n1840
* NET 3111 = abc_11867_new_n1839
* NET 3112 = abc_11867_new_n1838
* NET 3114 = abc_11867_new_n1826
* NET 3118 = abc_11867_new_n1861
* NET 3121 = abc_11867_new_n1886
* NET 3123 = abc_11867_new_n1859
* NET 3127 = abc_11867_new_n1851
* NET 3128 = abc_11867_new_n1863
* NET 3129 = abc_11867_new_n1867
* NET 3130 = abc_11867_new_n1879
* NET 3134 = abc_11867_new_n1842
* NET 3135 = abc_11867_new_n1845
* NET 3137 = abc_11867_new_n1710
* NET 3139 = abc_11867_new_n1870
* NET 3141 = abc_11867_new_n1871
* NET 3143 = abc_11867_new_n1872
* NET 3145 = abc_11867_new_n1873
* NET 3146 = abc_11867_new_n1869
* NET 3148 = abc_11867_new_n848
* NET 3150 = abc_11867_new_n503
* NET 3156 = abc_11867_new_n778
* NET 3158 = abc_11867_new_n588
* NET 3165 = abc_11867_new_n779
* NET 3167 = abc_11867_new_n772
* NET 3170 = abc_11867_new_n504
* NET 3171 = abc_11867_new_n510
* NET 3172 = abc_11867_new_n597
* NET 3175 = abc_11867_new_n428_hfns_5
* NET 3177 = abc_11867_new_n811
* NET 3179 = abc_11867_new_n485_hfns_4
* NET 3182 = abc_11867_new_n528
* NET 3184 = abc_11867_new_n737
* NET 3186 = abc_11867_new_n669
* NET 3187 = abc_11867_new_n554
* NET 3191 = abc_11867_new_n790
* NET 3192 = abc_11867_new_n781
* NET 3193 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[2]
* NET 3197 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[1]
* NET 3226 = subckt_1723_sff1_x4.y
* NET 3227 = subckt_1723_sff1_x4.sff_m
* NET 3229 = abc_11867_new_n1684
* NET 3241 = subckt_1685_sff1_x4.y
* NET 3242 = subckt_1685_sff1_x4.sff_m
* NET 3244 = abc_11867_new_n773
* NET 3250 = abc_11867_new_n511
* NET 3251 = abc_11867_new_n489
* NET 3252 = abc_11867_new_n502
* NET 3253 = abc_11867_new_n711
* NET 3258 = abc_11867_new_n839
* NET 3260 = abc_11867_new_n780
* NET 3261 = abc_11867_new_n529
* NET 3264 = abc_11867_new_n816
* NET 3267 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[0]
* NET 3268 = abc_11867_new_n815
* NET 3270 = subckt_1628_sff1_x4.y
* NET 3271 = subckt_1628_sff1_x4.sff_m
* NET 3275 = abc_11867_new_n1918
* NET 3276 = abc_11867_new_n1917
* NET 3279 = subckt_1723_sff1_x4.sff_s
* NET 3282 = abc_11867_auto_rtlil_cc_2608_muxgate_11794
* NET 3283 = subckt_1723_sff1_x4.ckr
* NET 3284 = subckt_1723_sff1_x4.u
* NET 3285 = subckt_1723_sff1_x4.nckr
* NET 3286 = abc_11867_new_n1790
* NET 3287 = abc_11867_new_n1901
* NET 3293 = abc_11867_new_n1733
* NET 3300 = a[6]
* NET 3303 = abc_11867_new_n1780
* NET 3307 = abc_11867_new_n1781
* NET 3310 = abc_11867_new_n1888
* NET 3313 = abc_11867_new_n1890
* NET 3315 = abc_11867_new_n1680
* NET 3316 = abc_11867_new_n1804
* NET 3320 = abc_11867_new_n1730
* NET 3327 = abc_11867_new_n1850
* NET 3330 = abc_11867_new_n1852
* NET 3340 = abc_11867_new_n1882
* NET 3348 = abc_11867_new_n1682
* NET 3353 = abc_11867_new_n1679
* NET 3356 = abc_11867_new_n1708
* NET 3361 = abc_11867_new_n1678
* NET 3370 = abc_11867_new_n636
* NET 3371 = abc_11867_new_n474
* NET 3373 = abc_11867_new_n520
* NET 3378 = abc_11867_new_n643
* NET 3379 = abc_11867_new_n637
* NET 3382 = subckt_1685_sff1_x4.sff_s
* NET 3384 = mos6502_src_reg[0]
* NET 3386 = subckt_1685_sff1_x4.u
* NET 3387 = subckt_1685_sff1_x4.ckr
* NET 3388 = subckt_1685_sff1_x4.nckr
* NET 3390 = abc_11867_new_n709
* NET 3391 = abc_11867_new_n386
* NET 3393 = abc_11867_new_n869
* NET 3399 = abc_11867_new_n596
* NET 3404 = abc_11867_new_n803
* NET 3405 = abc_11867_new_n807
* NET 3409 = abc_11867_new_n512
* NET 3410 = abc_11867_new_n513
* NET 3415 = abc_11867_new_n552
* NET 3416 = abc_11867_new_n553
* NET 3419 = abc_11867_new_n820
* NET 3421 = subckt_1628_sff1_x4.sff_s
* NET 3423 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[3]
* NET 3424 = subckt_1628_sff1_x4.ckr
* NET 3425 = subckt_1628_sff1_x4.u
* NET 3426 = subckt_1628_sff1_x4.nckr
* NET 3507 = abc_11867_new_n1549
* NET 3508 = abc_11867_auto_rtlil_cc_2608_muxgate_11828
* NET 3511 = abc_11867_auto_rtlil_cc_2608_muxgate_11826
* NET 3514 = subckt_1722_sff1_x4.sff_s
* NET 3515 = subckt_1722_sff1_x4.y
* NET 3517 = subckt_1722_sff1_x4.sff_m
* NET 3519 = abc_11867_auto_rtlil_cc_2608_muxgate_11792
* NET 3520 = subckt_1722_sff1_x4.u
* NET 3521 = subckt_1722_sff1_x4.ckr
* NET 3522 = subckt_1722_sff1_x4.nckr
* NET 3523 = subckt_1754_sff1_x4.sff_s
* NET 3525 = subckt_1754_sff1_x4.y
* NET 3526 = subckt_1754_sff1_x4.sff_m
* NET 3529 = subckt_1754_sff1_x4.u
* NET 3530 = subckt_1754_sff1_x4.nckr
* NET 3531 = subckt_1754_sff1_x4.ckr
* NET 3532 = abc_11867_new_n1140
* NET 3537 = abc_11867_new_n1146
* NET 3542 = abc_11867_new_n1686
* NET 3543 = abc_11867_new_n1787
* NET 3546 = abc_11867_new_n1806
* NET 3552 = abc_11867_new_n1712
* NET 3553 = abc_11867_new_n1715
* NET 3556 = abc_11867_new_n1650
* NET 3559 = abc_11867_new_n1805
* NET 3562 = abc_11867_new_n1797
* NET 3566 = abc_11867_new_n1731
* NET 3567 = abc_11867_new_n1857
* NET 3569 = abc_11867_new_n1858
* NET 3570 = abc_11867_new_n1860
* NET 3571 = abc_11867_new_n1849
* NET 3575 = abc_11867_new_n1885
* NET 3577 = abc_11867_new_n1887
* NET 3579 = abc_11867_new_n1701
* NET 3581 = abc_11867_new_n1702
* NET 3582 = abc_11867_new_n847
* NET 3583 = abc_11867_new_n845
* NET 3586 = abc_11867_new_n1709
* NET 3587 = abc_11867_new_n1707
* NET 3593 = subckt_1715_sff1_x4.sff_s
* NET 3595 = subckt_1715_sff1_x4.y
* NET 3596 = abc_11867_auto_rtlil_cc_2608_muxgate_11778
* NET 3598 = subckt_1715_sff1_x4.sff_m
* NET 3599 = subckt_1715_sff1_x4.nckr
* NET 3600 = subckt_1715_sff1_x4.u
* NET 3601 = subckt_1715_sff1_x4.ckr
* NET 3602 = abc_11867_new_n356
* NET 3603 = abc_11867_new_n1654
* NET 3606 = abc_11867_new_n1658
* NET 3608 = abc_11867_new_n765
* NET 3610 = abc_11867_new_n1647
* NET 3611 = abc_11867_new_n1653
* NET 3613 = abc_11867_new_n1652
* NET 3618 = abc_11867_new_n740
* NET 3622 = abc_11867_new_n866
* NET 3623 = abc_11867_new_n501
* NET 3624 = abc_11867_new_n713
* NET 3625 = abc_11867_new_n710
* NET 3628 = abc_11867_new_n712
* NET 3629 = abc_11867_new_n714
* NET 3635 = abc_11867_new_n703
* NET 3636 = abc_11867_new_n702
* NET 3639 = abc_11867_new_n589
* NET 3641 = abc_11867_new_n808
* NET 3642 = abc_11867_new_n826
* NET 3644 = abc_11867_new_n789
* NET 3645 = abc_11867_new_n788
* NET 3650 = abc_11867_new_n716
* NET 3651 = abc_11867_new_n715
* NET 3656 = abc_11867_new_n818
* NET 3659 = abc_11867_new_n819
* NET 3660 = abc_11867_new_n827
* NET 3661 = flatten_mos6502_auto_fsm_map_cc_288_map_fsm_1405_y[4]
* NET 3662 = abc_11867_new_n478
* NET 3664 = abc_11867_new_n814
* NET 3665 = abc_11867_new_n792
* NET 3667 = abc_11867_new_n802
* NET 3701 = subckt_1759_sff1_x4.sff_s
* NET 3703 = subckt_1759_sff1_x4.y
* NET 3705 = subckt_1759_sff1_x4.sff_m
* NET 3707 = subckt_1759_sff1_x4.u
* NET 3708 = clk_root_tr_0
* NET 3709 = subckt_1759_sff1_x4.nckr
* NET 3710 = subckt_1759_sff1_x4.ckr
* NET 3711 = abc_11867_new_n1036
* NET 3714 = abc_11867_new_n1031
* NET 3716 = abc_11867_new_n355
* NET 3717 = abc_11867_new_n1932
* NET 3718 = abc_11867_auto_rtlil_cc_2608_muxgate_11856
* NET 3720 = abc_11867_new_n1900
* NET 3722 = abc_11867_new_n1933
* NET 3723 = abc_11867_new_n1023
* NET 3725 = abc_11867_new_n1752
* NET 3730 = abc_11867_new_n1753
* NET 3735 = abc_11867_new_n1755
* NET 3737 = abc_11867_new_n1711
* NET 3740 = abc_11867_new_n1809
* NET 3743 = abc_11867_new_n1810
* NET 3744 = abc_11867_new_n1714
* NET 3748 = abc_11867_new_n1801
* NET 3750 = abc_11867_new_n1921
* NET 3751 = abc_11867_new_n1919
* NET 3752 = abc_11867_new_n1922
* NET 3754 = abc_11867_new_n1803
* NET 3757 = abc_11867_new_n1774
* NET 3759 = abc_11867_new_n1824
* NET 3763 = abc_11867_new_n1848
* NET 3765 = abc_11867_new_n1539
* NET 3768 = abc_11867_new_n1865
* NET 3771 = abc_11867_new_n968
* NET 3774 = abc_11867_new_n1703
* NET 3776 = abc_11867_new_n841
* NET 3780 = abc_11867_new_n1648
* NET 3782 = abc_11867_new_n1704
* NET 3783 = abc_11867_new_n1706
* NET 3787 = mos6502_backwards
* NET 3788 = abc_11867_new_n1705
* NET 3792 = reset
* NET 3794 = abc_11867_new_n846
* NET 3797 = abc_11867_new_n974
* NET 3801 = abc_11867_new_n969
* NET 3802 = abc_11867_new_n1657
* NET 3804 = abc_11867_new_n1655
* NET 3809 = abc_11867_new_n564
* NET 3812 = abc_11867_new_n624
* NET 3819 = abc_11867_new_n1651
* NET 3826 = abc_11867_new_n494
* NET 3828 = subckt_1684_sff1_x4.sff_s
* NET 3829 = subckt_1684_sff1_x4.y
* NET 3831 = subckt_1684_sff1_x4.sff_m
* NET 3832 = subckt_1684_sff1_x4.u
* NET 3834 = clk_root_tl_0
* NET 3835 = subckt_1684_sff1_x4.ckr
* NET 3836 = subckt_1684_sff1_x4.nckr
* NET 3839 = abc_11867_new_n497
* NET 3841 = abc_11867_new_n784
* NET 3842 = abc_11867_new_n568
* NET 3844 = abc_11867_new_n594
* NET 3847 = abc_11867_new_n692
* NET 3850 = abc_11867_new_n693
* NET 3851 = abc_11867_new_n694
* NET 3853 = abc_11867_new_n787
* NET 3856 = abc_11867_new_n739
* NET 3857 = abc_11867_new_n426_hfns_0
* NET 3858 = abc_11867_new_n762
* NET 3860 = abc_11867_new_n732
* NET 3863 = abc_11867_new_n731
* NET 3865 = abc_11867_new_n838
* NET 3867 = abc_11867_new_n785
* NET 3868 = abc_11867_new_n786
* NET 3871 = abc_11867_new_n813
* NET 3872 = abc_11867_new_n812
* NET 3876 = abc_11867_new_n801
* NET 3877 = abc_11867_new_n799
* NET 3955 = abc_11867_auto_rtlil_cc_2608_muxgate_11866
* NET 3956 = mos6502_alu_ai7
* NET 3958 = abc_11867_new_n1677
* NET 3962 = abc_11867_auto_rtlil_cc_2608_muxgate_11858
* NET 3964 = abc_11867_new_n1916
* NET 3968 = abc_11867_new_n1136
* NET 3969 = abc_11867_new_n1020
* NET 3971 = abc_11867_new_n1931
* NET 3972 = abc_11867_new_n1015
* NET 3978 = abc_11867_new_n1132
* NET 3986 = abc_11867_new_n1807
* NET 3987 = abc_11867_new_n1777
* NET 3989 = abc_11867_new_n1778
* NET 3990 = abc_11867_new_n1776
* NET 3991 = abc_11867_new_n1800
* NET 3993 = abc_11867_new_n1775
* NET 3995 = abc_11867_new_n1773
* NET 3997 = abc_11867_new_n1769
* NET 3999 = abc_11867_new_n1110
* NET 4003 = abc_11867_new_n1819
* NET 4007 = abc_11867_new_n1868
* NET 4009 = abc_11867_new_n353
* NET 4012 = abc_11867_new_n1126
* NET 4018 = abc_11867_new_n1043
* NET 4021 = abc_11867_new_n727
* NET 4022 = clk
* NET 4024 = abc_11867_new_n849
* NET 4025 = abc_11867_new_n918
* NET 4029 = abc_11867_new_n919
* NET 4030 = abc_11867_new_n357
* NET 4032 = abc_11867_new_n347
* NET 4033 = abc_11867_new_n1656
* NET 4036 = subckt_1675_sff1_x4.sff_s
* NET 4037 = subckt_1675_sff1_x4.y
* NET 4039 = subckt_1675_sff1_x4.sff_m
* NET 4041 = subckt_1675_sff1_x4.u
* NET 4042 = subckt_1675_sff1_x4.ckr
* NET 4043 = subckt_1675_sff1_x4.nckr
* NET 4045 = abc_11867_new_n514
* NET 4047 = abc_11867_new_n496
* NET 4048 = abc_11867_new_n498
* NET 4049 = abc_11867_new_n514_hfns_2
* NET 4051 = abc_11867_new_n485_hfns_3
* NET 4054 = subckt_1687_sff1_x4.sff_s
* NET 4055 = subckt_1687_sff1_x4.y
* NET 4058 = subckt_1687_sff1_x4.sff_m
* NET 4059 = subckt_1687_sff1_x4.u
* NET 4060 = subckt_1687_sff1_x4.ckr
* NET 4061 = abc_11867_new_n492
* NET 4062 = subckt_1687_sff1_x4.nckr
* NET 4067 = abc_11867_new_n471_hfns_1
* NET 4068 = abc_11867_new_n482_hfns_0
* NET 4070 = abc_11867_new_n704
* NET 4071 = abc_11867_new_n699
* NET 4074 = abc_11867_new_n822
* NET 4075 = abc_11867_new_n426_hfns_1
* NET 4076 = abc_11867_new_n478_hfns_3
* NET 4078 = abc_11867_new_n683
* NET 4079 = rdy
* NET 4120 = subckt_1741_sff1_x4.sff_s
* NET 4122 = subckt_1741_sff1_x4.y
* NET 4124 = subckt_1741_sff1_x4.sff_m
* NET 4125 = subckt_1741_sff1_x4.u
* NET 4127 = subckt_1741_sff1_x4.ckr
* NET 4128 = subckt_1741_sff1_x4.nckr
* NET 4129 = abc_11867_new_n1032
* NET 4130 = abc_11867_new_n1035
* NET 4133 = abc_11867_new_n1034
* NET 4134 = abc_11867_new_n375
* NET 4137 = abc_11867_new_n1005
* NET 4141 = abc_11867_new_n1808
* NET 4143 = abc_11867_new_n1811
* NET 4149 = abc_11867_new_n1815
* NET 4152 = abc_11867_new_n1893
* NET 4155 = abc_11867_new_n1812
* NET 4156 = abc_11867_new_n1898
* NET 4157 = abc_11867_new_n1813
* NET 4160 = abc_11867_new_n1124
* NET 4166 = abc_11867_new_n1823
* NET 4167 = abc_11867_new_n473_hfns_2
* NET 4171 = abc_11867_new_n1795
* NET 4172 = abc_11867_new_n1416
* NET 4173 = abc_11867_new_n1690
* NET 4176 = abc_11867_new_n1118
* NET 4178 = abc_11867_new_n610
* NET 4183 = abc_11867_new_n1820
* NET 4184 = abc_11867_new_n997
* NET 4186 = abc_11867_new_n928
* NET 4189 = abc_11867_new_n1866
* NET 4191 = abc_11867_new_n933
* NET 4192 = abc_11867_new_n931
* NET 4193 = abc_11867_new_n932
* NET 4197 = abc_11867_new_n968_hfns_2
* NET 4198 = abc_11867_new_n1012
* NET 4202 = abc_11867_new_n920
* NET 4203 = abc_11867_new_n843
* NET 4206 = abc_11867_new_n921
* NET 4207 = abc_11867_new_n924
* NET 4208 = abc_11867_new_n923
* NET 4212 = abc_11867_new_n922
* NET 4224 = abc_11867_new_n1497
* NET 4228 = abc_11867_new_n728
* NET 4230 = irq
* NET 4234 = abc_11867_new_n1392
* NET 4236 = abc_11867_new_n1337
* NET 4241 = subckt_1709_sff1_x4.sff_s
* NET 4242 = subckt_1709_sff1_x4.y
* NET 4244 = abc_11867_auto_rtlil_cc_2608_muxgate_11768
* NET 4245 = subckt_1709_sff1_x4.sff_m
* NET 4247 = subckt_1709_sff1_x4.u
* NET 4248 = subckt_1709_sff1_x4.ckr
* NET 4249 = subckt_1709_sff1_x4.nckr
* NET 4251 = abc_11867_new_n385
* NET 4254 = abc_11867_auto_rtlil_cc_2608_muxgate_11708
* NET 4255 = mos6502_shift_right
* NET 4260 = abc_11867_new_n346
* NET 4262 = subckt_1680_sff1_x4.sff_s
* NET 4263 = subckt_1680_sff1_x4.y
* NET 4266 = subckt_1680_sff1_x4.sff_m
* NET 4267 = subckt_1680_sff1_x4.ckr
* NET 4268 = subckt_1680_sff1_x4.u
* NET 4269 = subckt_1680_sff1_x4.nckr
* NET 4270 = mos6502_index_y
* NET 4271 = abc_11867_auto_rtlil_cc_2608_muxgate_11728
* NET 4276 = abc_11867_new_n805
* NET 4280 = abc_11867_new_n783
* NET 4286 = abc_11867_new_n684
* NET 4287 = abc_11867_new_n686
* NET 4292 = abc_11867_new_n782
* NET 4293 = abc_11867_new_n475_hfns_0
* NET 4295 = abc_11867_new_n514_hfns_0
* NET 4298 = abc_11867_new_n717
* NET 4299 = abc_11867_new_n720
* NET 4302 = abc_11867_new_n475_hfns_1
* NET 4306 = abc_11867_new_n471_hfns_0
* NET 4310 = abc_11867_new_n608_hfns_0
* NET 4311 = abc_11867_new_n548
* NET 4312 = abc_11867_new_n531
* NET 4315 = abc_11867_new_n796
* NET 4317 = abc_11867_new_n794
* NET 4318 = abc_11867_new_n795
* NET 4402 = abc_11867_new_n1134
* NET 4403 = abc_11867_new_n1139
* NET 4405 = abc_11867_new_n1000
* NET 4406 = abc_11867_new_n351
* NET 4413 = abc_11867_new_n354
* NET 4414 = abc_11867_new_n1123
* NET 4416 = abc_11867_new_n1897
* NET 4418 = abc_11867_new_n1033
* NET 4424 = abc_11867_new_n1847
* NET 4426 = abc_11867_new_n1802
* NET 4427 = abc_11867_new_n891
* NET 4428 = abc_11867_new_n992
* NET 4429 = abc_11867_new_n954_hfns_1
* NET 4433 = abc_11867_new_n1038
* NET 4437 = abc_11867_new_n905
* NET 4438 = abc_11867_new_n930
* NET 4439 = abc_11867_new_n1007
* NET 4447 = abc_11867_new_n1399
* NET 4448 = abc_11867_new_n1366
* NET 4449 = abc_11867_new_n1368
* NET 4460 = abc_11867_auto_rtlil_cc_2608_muxgate_11734
* NET 4461 = mos6502_dst_reg[0]
* NET 4468 = abc_11867_new_n630
* NET 4470 = abc_11867_new_n633
* NET 4472 = abc_11867_new_n679
* NET 4473 = abc_11867_new_n719
* NET 4474 = abc_11867_new_n682
* NET 4476 = abc_11867_new_n723
* NET 4477 = abc_11867_new_n678
* NET 4479 = abc_11867_new_n793
* NET 4480 = subckt_1745_sff1_x4.sff_s
* NET 4481 = subckt_1745_sff1_x4.y
* NET 4482 = subckt_1745_sff1_x4.sff_m
* NET 4483 = subckt_1745_sff1_x4.u
* NET 4484 = subckt_1745_sff1_x4.ckr
* NET 4485 = subckt_1745_sff1_x4.nckr
* NET 4489 = abc_11867_new_n1138
* NET 4491 = subckt_1615_nmx2_x1.q
* NET 4492 = abc_11867_new_n1899
* NET 4497 = abc_11867_new_n1814
* NET 4498 = abc_11867_new_n1891
* NET 4502 = abc_11867_new_n1895
* NET 4503 = abc_11867_new_n1894
* NET 4507 = abc_11867_new_n423
* NET 4510 = abc_11867_new_n1681
* NET 4511 = abc_11867_new_n1799
* NET 4512 = abc_11867_new_n1798
* NET 4517 = abc_11867_new_n647
* NET 4518 = abc_11867_new_n609
* NET 4525 = abc_11867_new_n619
* NET 4527 = abc_11867_new_n577
* NET 4529 = abc_11867_new_n1471
* NET 4530 = abc_11867_new_n434
* NET 4531 = subckt_1689_sff1_x4.sff_s
* NET 4532 = subckt_1689_sff1_x4.ckr
* NET 4533 = subckt_1689_sff1_x4.y
* NET 4534 = subckt_1689_sff1_x4.sff_m
* NET 4535 = subckt_1689_sff1_x4.u
* NET 4536 = subckt_1689_sff1_x4.nckr
* NET 4537 = abc_11867_new_n1404
* NET 4538 = mos6502_nmi_edge
* NET 4540 = abc_11867_new_n617
* NET 4542 = subckt_1672_sff1_x4.sff_s
* NET 4543 = mos6502_op[2]
* NET 4544 = subckt_1672_sff1_x4.y
* NET 4545 = subckt_1672_sff1_x4.sff_m
* NET 4546 = subckt_1672_sff1_x4.u
* NET 4547 = subckt_1672_sff1_x4.ckr
* NET 4548 = abc_11867_new_n587
* NET 4549 = subckt_1672_sff1_x4.nckr
* NET 4552 = abc_11867_new_n1181
* NET 4556 = abc_11867_new_n358
* NET 4557 = subckt_1686_sff1_x4.sff_s
* NET 4558 = mos6502_src_reg[1]
* NET 4559 = subckt_1686_sff1_x4.y
* NET 4560 = subckt_1686_sff1_x4.sff_m
* NET 4561 = subckt_1686_sff1_x4.u
* NET 4562 = subckt_1686_sff1_x4.ckr
* NET 4563 = subckt_1686_sff1_x4.nckr
* NET 4564 = subckt_1682_sff1_x4.sff_s
* NET 4565 = subckt_1682_sff1_x4.sff_m
* NET 4566 = subckt_1682_sff1_x4.u
* NET 4567 = subckt_1682_sff1_x4.ckr
* NET 4568 = subckt_1682_sff1_x4.y
* NET 4569 = subckt_1682_sff1_x4.nckr
* NET 4570 = abc_11867_auto_rtlil_cc_2608_muxgate_11724
* NET 4572 = abc_11867_new_n475_hfns_2
* NET 4573 = abc_11867_new_n482_hfns_1
* NET 4574 = abc_11867_new_n473_hfns_0
* NET 4575 = abc_11867_new_n514_hfns_1
* NET 4577 = abc_11867_new_n626
* NET 4579 = abc_11867_new_n680
* NET 4582 = abc_11867_new_n671
* NET 4583 = abc_11867_new_n533
* NET 4612 = subckt_1758_sff1_x4.y
* NET 4614 = subckt_1758_sff1_x4.sff_m
* NET 4615 = subckt_1758_sff1_x4.ckr
* NET 4617 = subckt_1751_sff1_x4.y
* NET 4619 = subckt_1751_sff1_x4.sff_m
* NET 4620 = subckt_1751_sff1_x4.ckr
* NET 4624 = subckt_1697_sff1_x4.y
* NET 4626 = subckt_1697_sff1_x4.sff_m
* NET 4627 = subckt_1697_sff1_x4.ckr
* NET 4631 = subckt_1674_sff1_x4.y
* NET 4633 = subckt_1674_sff1_x4.sff_m
* NET 4634 = subckt_1674_sff1_x4.ckr
* NET 4635 = abc_11867_new_n387
* NET 4641 = abc_11867_auto_rtlil_cc_2608_muxgate_11862
* NET 4644 = abc_11867_new_n1915
* NET 4647 = abc_11867_new_n1016
* NET 4648 = abc_11867_new_n1019
* NET 4651 = abc_11867_new_n1130
* NET 4658 = abc_11867_new_n1142
* NET 4662 = abc_11867_new_n1145
* NET 4663 = abc_11867_new_n1144
* NET 4665 = subckt_1758_sff1_x4.sff_s
* NET 4666 = abc_11867_auto_rtlil_cc_2608_muxgate_11864
* NET 4668 = subckt_1758_sff1_x4.u
* NET 4669 = subckt_1758_sff1_x4.nckr
* NET 4672 = abc_11867_new_n1122
* NET 4680 = subckt_1751_sff1_x4.sff_s
* NET 4681 = abc_11867_auto_rtlil_cc_2608_muxgate_11850
* NET 4683 = subckt_1751_sff1_x4.nckr
* NET 4684 = subckt_1751_sff1_x4.u
* NET 4685 = abc_11867_new_n1794
* NET 4688 = abc_11867_new_n1772
* NET 4690 = abc_11867_new_n1771
* NET 4693 = abc_11867_new_n981
* NET 4698 = abc_11867_new_n1109
* NET 4701 = abc_11867_new_n422
* NET 4702 = subckt_1697_sff1_x4.sff_s
* NET 4704 = subckt_1697_sff1_x4.u
* NET 4705 = abc_11867_new_n352
* NET 4706 = subckt_1697_sff1_x4.nckr
* NET 4707 = abc_11867_new_n1474
* NET 4712 = di[7]
* NET 4714 = mos6502_dihold[7]
* NET 4715 = subckt_101_nmx2_x1.q
* NET 4717 = abc_11867_new_n1488
* NET 4720 = mos6502_res
* NET 4721 = abc_11867_auto_rtlil_cc_2608_muxgate_11740
* NET 4722 = abc_11867_new_n323
* NET 4725 = abc_11867_new_n1393
* NET 4727 = abc_11867_new_n1401
* NET 4728 = abc_11867_new_n1400
* NET 4730 = abc_11867_new_n363
* NET 4731 = abc_11867_new_n324
* NET 4734 = mos6502_write_back
* NET 4735 = abc_11867_new_n1394
* NET 4737 = abc_11867_new_n1339
* NET 4738 = abc_11867_new_n1338
* NET 4739 = abc_11867_new_n331
* NET 4742 = abc_11867_new_n328
* NET 4744 = abc_11867_new_n1398
* NET 4749 = abc_11867_new_n1365
* NET 4752 = subckt_1674_sff1_x4.sff_s
* NET 4754 = subckt_1674_sff1_x4.u
* NET 4755 = subckt_1674_sff1_x4.nckr
* NET 4756 = abc_11867_new_n1298
* NET 4757 = abc_11867_auto_rtlil_cc_2608_muxgate_11730
* NET 4759 = abc_11867_auto_rtlil_cc_2608_muxgate_11706
* NET 4760 = mos6502_rotate
* NET 4765 = abc_11867_auto_rtlil_cc_2608_muxgate_11732
* NET 4766 = abc_11867_new_n1300
* NET 4769 = abc_11867_auto_rtlil_cc_2608_muxgate_11720
* NET 4770 = mos6502_inc
* NET 4779 = abc_11867_new_n470
* NET 4782 = abc_11867_new_n458
* NET 4786 = abc_11867_new_n457
* NET 4788 = abc_11867_new_n1291
* NET 4790 = abc_11867_new_n532
* NET 4792 = abc_11867_new_n688
* NET 4795 = abc_11867_new_n718
* NET 4798 = abc_11867_new_n761
* NET 4801 = abc_11867_new_n746
* NET 4802 = abc_11867_new_n722
* NET 4803 = abc_11867_new_n744
* NET 4885 = abc_11867_new_n1547
* NET 4887 = subckt_1753_sff1_x4.sff_s
* NET 4888 = subckt_1753_sff1_x4.y
* NET 4890 = subckt_1753_sff1_x4.sff_m
* NET 4892 = subckt_1753_sff1_x4.u
* NET 4893 = subckt_1753_sff1_x4.ckr
* NET 4894 = subckt_1753_sff1_x4.nckr
* NET 4895 = abc_11867_new_n1143
* NET 4896 = abc_11867_new_n341
* NET 4898 = abc_11867_new_n1004
* NET 4900 = abc_11867_new_n1121
* NET 4901 = abc_11867_new_n336
* NET 4902 = abc_11867_new_n335
* NET 4905 = subckt_1752_sff1_x4.sff_s
* NET 4906 = subckt_1752_sff1_x4.y
* NET 4909 = subckt_1752_sff1_x4.sff_m
* NET 4910 = subckt_1752_sff1_x4.u
* NET 4911 = subckt_1752_sff1_x4.ckr
* NET 4912 = subckt_1752_sff1_x4.nckr
* NET 4913 = abc_11867_auto_rtlil_cc_2608_muxgate_11852
* NET 4914 = abc_11867_new_n1896
* NET 4921 = abc_11867_new_n1112
* NET 4924 = abc_11867_new_n1116
* NET 4925 = abc_11867_new_n1117
* NET 4927 = abc_11867_new_n944
* NET 4929 = do[7]
* NET 4932 = abc_11867_new_n890
* NET 4934 = abc_11867_new_n976
* NET 4939 = abc_11867_new_n333
* NET 4942 = abc_11867_new_n929
* NET 4945 = abc_11867_new_n887
* NET 4947 = abc_11867_new_n1844
* NET 4951 = abc_11867_new_n619_hfns_2
* NET 4953 = abc_11867_new_n888
* NET 4955 = mos6502_i
* NET 4956 = abc_11867_new_n903
* NET 4958 = subckt_1713_sff1_x4.sff_s
* NET 4960 = subckt_1713_sff1_x4.y
* NET 4961 = subckt_1713_sff1_x4.sff_m
* NET 4963 = abc_11867_auto_rtlil_cc_2608_muxgate_11776
* NET 4965 = subckt_1713_sff1_x4.u
* NET 4966 = subckt_1713_sff1_x4.nckr
* NET 4967 = subckt_1713_sff1_x4.ckr
* NET 4969 = subckt_1670_sff1_x4.sff_s
* NET 4970 = subckt_1670_sff1_x4.y
* NET 4973 = subckt_1670_sff1_x4.sff_m
* NET 4974 = subckt_1670_sff1_x4.u
* NET 4975 = subckt_1670_sff1_x4.ckr
* NET 4976 = subckt_1670_sff1_x4.nckr
* NET 4978 = subckt_1699_sff1_x4.sff_s
* NET 4979 = subckt_1699_sff1_x4.y
* NET 4982 = subckt_1699_sff1_x4.sff_m
* NET 4983 = abc_11867_auto_rtlil_cc_2608_muxgate_11746
* NET 4984 = subckt_1699_sff1_x4.u
* NET 4985 = subckt_1699_sff1_x4.ckr
* NET 4986 = subckt_1699_sff1_x4.nckr
* NET 4987 = abc_11867_new_n1367
* NET 4995 = abc_11867_new_n1181_hfns_2
* NET 4997 = abc_11867_new_n764
* NET 4998 = abc_11867_new_n1363
* NET 4999 = abc_11867_new_n344
* NET 5000 = abc_11867_new_n384
* NET 5002 = abc_11867_new_n1297
* NET 5003 = mos6502_php
* NET 5005 = subckt_1661_sff1_x4.sff_s
* NET 5006 = subckt_1661_sff1_x4.y
* NET 5009 = subckt_1661_sff1_x4.sff_m
* NET 5010 = subckt_1661_sff1_x4.u
* NET 5011 = subckt_1661_sff1_x4.ckr
* NET 5012 = subckt_1661_sff1_x4.nckr
* NET 5013 = abc_11867_new_n1221
* NET 5015 = mos6502_dst_reg[1]
* NET 5017 = subckt_1688_sff1_x4.sff_s
* NET 5018 = subckt_1688_sff1_x4.y
* NET 5021 = subckt_1688_sff1_x4.sff_m
* NET 5022 = subckt_1688_sff1_x4.u
* NET 5023 = subckt_1688_sff1_x4.ckr
* NET 5024 = subckt_1688_sff1_x4.nckr
* NET 5025 = abc_11867_new_n388
* NET 5026 = abc_11867_new_n1317
* NET 5027 = abc_11867_auto_rtlil_cc_2608_muxgate_11736
* NET 5030 = abc_11867_new_n1315
* NET 5031 = abc_11867_new_n685
* NET 5032 = abc_11867_new_n697
* NET 5034 = abc_11867_new_n760
* NET 5036 = abc_11867_new_n748
* NET 5037 = abc_11867_new_n681
* NET 5038 = abc_11867_new_n677
* NET 5040 = abc_11867_new_n759
* NET 5041 = abc_11867_new_n756
* NET 5042 = abc_11867_new_n687
* NET 5044 = abc_11867_new_n628
* NET 5077 = abc_11867_new_n1559
* NET 5078 = abc_11867_new_n1546
* NET 5089 = abc_11867_new_n1001
* NET 5090 = abc_11867_auto_rtlil_cc_2608_muxgate_11854
* NET 5092 = abc_11867_new_n1892
* NET 5099 = abc_11867_new_n1675
* NET 5108 = mos6502_alu_hc
* NET 5109 = abc_11867_new_n1120
* NET 5110 = abc_11867_new_n1114
* NET 5113 = abc_11867_new_n1115
* NET 5114 = abc_11867_new_n1113
* NET 5118 = abc_11867_new_n1108
* NET 5120 = abc_11867_new_n1107
* NET 5121 = abc_11867_new_n1106
* NET 5124 = abc_11867_new_n1674
* NET 5129 = abc_11867_new_n372
* NET 5132 = abc_11867_new_n977
* NET 5133 = abc_11867_new_n980
* NET 5136 = abc_11867_new_n989
* NET 5139 = abc_11867_new_n985
* NET 5140 = abc_11867_new_n988
* NET 5143 = mos6502_abl[0]
* NET 5144 = abc_11867_new_n1481
* NET 5147 = abc_11867_new_n648
* NET 5148 = abc_11867_new_n611
* NET 5150 = abc_11867_new_n1011
* NET 5151 = abc_11867_new_n1010
* NET 5154 = abc_11867_new_n1008
* NET 5160 = abc_11867_new_n1496
* NET 5161 = abc_11867_new_n1498
* NET 5162 = abc_11867_new_n1499
* NET 5164 = abc_11867_new_n1673
* NET 5168 = abc_11867_new_n595
* NET 5169 = abc_11867_new_n631
* NET 5176 = abc_11867_new_n1099
* NET 5178 = abc_11867_new_n329
* NET 5180 = mos6502_op[0]
* NET 5181 = abc_11867_auto_rtlil_cc_2608_muxgate_11698
* NET 5186 = subckt_1673_sff1_x4.sff_s
* NET 5188 = rdy_hfns_4
* NET 5189 = subckt_1673_sff1_x4.y
* NET 5191 = subckt_1673_sff1_x4.sff_m
* NET 5193 = subckt_1673_sff1_x4.u
* NET 5194 = subckt_1673_sff1_x4.nckr
* NET 5195 = subckt_1673_sff1_x4.ckr
* NET 5196 = abc_11867_auto_rtlil_cc_2608_muxgate_11704
* NET 5197 = mos6502_op[3]
* NET 5202 = mos6502_cli
* NET 5204 = subckt_1666_sff1_x4.sff_s
* NET 5205 = subckt_1666_sff1_x4.y
* NET 5207 = subckt_1666_sff1_x4.sff_m
* NET 5209 = subckt_1666_sff1_x4.u
* NET 5210 = subckt_1666_sff1_x4.ckr
* NET 5211 = subckt_1666_sff1_x4.nckr
* NET 5212 = abc_11867_new_n1237
* NET 5213 = abc_11867_auto_rtlil_cc_2608_muxgate_11702
* NET 5216 = subckt_1667_sff1_x4.sff_s
* NET 5217 = subckt_1667_sff1_x4.y
* NET 5219 = subckt_1667_sff1_x4.sff_m
* NET 5221 = subckt_1667_sff1_x4.ckr
* NET 5222 = subckt_1667_sff1_x4.u
* NET 5223 = abc_11867_new_n1185
* NET 5224 = subckt_1667_sff1_x4.nckr
* NET 5226 = abc_11867_auto_rtlil_cc_2608_muxgate_11680
* NET 5227 = mos6502_load_only
* NET 5229 = subckt_1681_sff1_x4.sff_s
* NET 5230 = subckt_1681_sff1_x4.y
* NET 5232 = abc_11867_auto_rtlil_cc_2608_muxgate_11722
* NET 5234 = subckt_1681_sff1_x4.sff_m
* NET 5235 = subckt_1681_sff1_x4.ckr
* NET 5236 = subckt_1681_sff1_x4.u
* NET 5237 = subckt_1681_sff1_x4.nckr
* NET 5238 = abc_11867_new_n757
* NET 5241 = abc_11867_new_n1278
* NET 5242 = abc_11867_new_n1314
* NET 5245 = abc_11867_new_n629
* NET 5249 = abc_11867_new_n1313
* NET 5256 = abc_11867_new_n750
* NET 5262 = abc_11867_new_n459
* NET 5265 = abc_11867_new_n547
* NET 5269 = abc_11867_new_n698
* NET 5273 = abc_11867_new_n758
* NET 5372 = abc_11867_new_n1025
* NET 5373 = abc_11867_new_n419
* NET 5377 = abc_11867_new_n1137
* NET 5379 = abc_11867_new_n1018
* NET 5380 = abc_11867_new_n373
* NET 5383 = abc_11867_new_n1135
* NET 5384 = abc_11867_new_n1128
* NET 5387 = mos6502_abl[6]
* NET 5388 = abc_11867_new_n1531
* NET 5390 = abc_11867_new_n1129
* NET 5391 = abc_11867_new_n1131
* NET 5394 = mos6502_abl[5]
* NET 5395 = abc_11867_new_n1727
* NET 5399 = abc_11867_new_n904
* NET 5401 = abc_11867_new_n1749
* NET 5406 = abc_11867_new_n1671
* NET 5408 = abc_11867_new_n984
* NET 5413 = abc_11867_new_n349
* NET 5414 = abc_11867_new_n1491
* NET 5416 = abc_11867_new_n1500
* NET 5417 = abc_11867_new_n350
* NET 5419 = mos6502_abl[4]
* NET 5420 = abc_11867_new_n979
* NET 5421 = abc_11867_new_n368
* NET 5424 = abc_11867_new_n1480
* NET 5426 = abc_11867_new_n1461
* NET 5428 = abc_11867_new_n1482
* NET 5429 = abc_11867_new_n348
* NET 5432 = abc_11867_new_n1478
* NET 5434 = abc_11867_new_n585
* NET 5435 = mos6502_abl[2]
* NET 5436 = abc_11867_new_n1490
* NET 5437 = abc_11867_new_n1489
* NET 5440 = abc_11867_new_n987
* NET 5443 = mos6502_abl[1]
* NET 5444 = abc_11867_new_n369
* NET 5445 = abc_11867_new_n1098
* NET 5447 = abc_11867_new_n431_hfns_1
* NET 5449 = abc_11867_new_n1403
* NET 5453 = mos6502_alu_co
* NET 5459 = subckt_1671_sff1_x4.sff_s
* NET 5460 = subckt_1671_sff1_x4.y
* NET 5463 = subckt_1671_sff1_x4.sff_m
* NET 5464 = subckt_1671_sff1_x4.u
* NET 5465 = subckt_1671_sff1_x4.ckr
* NET 5466 = subckt_1671_sff1_x4.nckr
* NET 5467 = abc_11867_new_n1397
* NET 5470 = subckt_1676_sff1_x4.sff_s
* NET 5471 = subckt_1676_sff1_x4.y
* NET 5474 = subckt_1676_sff1_x4.sff_m
* NET 5475 = subckt_1676_sff1_x4.u
* NET 5476 = subckt_1676_sff1_x4.nckr
* NET 5477 = subckt_1676_sff1_x4.ckr
* NET 5478 = abc_11867_auto_rtlil_cc_2608_muxgate_11710
* NET 5483 = abc_11867_new_n430_hfns_0
* NET 5485 = mos6502_sei
* NET 5486 = abc_11867_new_n1204
* NET 5487 = abc_11867_auto_rtlil_cc_2608_muxgate_11690
* NET 5489 = abc_11867_new_n1207
* NET 5490 = abc_11867_auto_rtlil_cc_2608_muxgate_11692
* NET 5492 = abc_11867_new_n557
* NET 5494 = abc_11867_new_n1205
* NET 5495 = abc_11867_new_n1257
* NET 5496 = abc_11867_new_n559
* NET 5498 = abc_11867_new_n1256
* NET 5500 = abc_11867_new_n1305
* NET 5501 = abc_11867_new_n1306
* NET 5502 = abc_11867_new_n1277
* NET 5503 = abc_11867_new_n1239
* NET 5504 = abc_11867_new_n1320
* NET 5505 = abc_11867_new_n749
* NET 5507 = abc_11867_new_n1319
* NET 5508 = abc_11867_new_n1318
* NET 5509 = abc_11867_new_n747
* NET 5551 = abc_11867_new_n418
* NET 5553 = abc_11867_new_n1532
* NET 5558 = abc_11867_new_n1358
* NET 5562 = abc_11867_new_n1540
* NET 5563 = mos6502_abl[7]
* NET 5566 = abc_11867_new_n1003
* NET 5567 = abc_11867_new_n371
* NET 5571 = mos6502_abl[3]
* NET 5574 = abc_11867_new_n619_hfns_1
* NET 5576 = abc_11867_new_n1506
* NET 5579 = subckt_1733_sff1_x4.sff_s
* NET 5580 = subckt_1733_sff1_x4.y
* NET 5582 = subckt_1733_sff1_x4.sff_m
* NET 5583 = subckt_1733_sff1_x4.u
* NET 5585 = subckt_1733_sff1_x4.ckr
* NET 5586 = subckt_1733_sff1_x4.nckr
* NET 5587 = abc_11867_new_n1487
* NET 5588 = abc_11867_new_n1493
* NET 5589 = abc_11867_auto_rtlil_cc_2608_muxgate_11814
* NET 5592 = subckt_1732_sff1_x4.sff_s
* NET 5593 = subckt_1732_sff1_x4.y
* NET 5594 = subckt_1732_sff1_x4.sff_m
* NET 5597 = subckt_1732_sff1_x4.ckr
* NET 5598 = subckt_1732_sff1_x4.u
* NET 5599 = subckt_1732_sff1_x4.nckr
* NET 5600 = abc_11867_new_n947
* NET 5603 = mos6502_pc[0]
* NET 5606 = mos6502_adj_bcd
* NET 5608 = subckt_1714_sff1_x4.sff_s
* NET 5609 = subckt_1714_sff1_x4.y
* NET 5612 = subckt_1714_sff1_x4.sff_m
* NET 5613 = subckt_1714_sff1_x4.ckr
* NET 5614 = subckt_1714_sff1_x4.u
* NET 5615 = subckt_1714_sff1_x4.nckr
* NET 5616 = abc_11867_new_n1484
* NET 5618 = abc_11867_new_n1464
* NET 5619 = abc_11867_new_n1470
* NET 5620 = abc_11867_new_n1469
* NET 5624 = abc_11867_new_n471_hfns_2
* NET 5628 = abc_11867_new_n1476
* NET 5629 = abc_11867_new_n1463
* NET 5632 = abc_11867_new_n370
* NET 5633 = abc_11867_new_n973
* NET 5637 = abc_11867_new_n1351
* NET 5641 = abc_11867_new_n879
* NET 5642 = abc_11867_new_n1375
* NET 5644 = abc_11867_new_n1378
* NET 5648 = abc_11867_new_n473_hfns_1
* NET 5653 = abc_11867_new_n376
* NET 5654 = abc_11867_new_n431_hfns_0
* NET 5658 = abc_11867_new_n1402
* NET 5664 = mos6502_compare
* NET 5665 = abc_11867_new_n1395
* NET 5668 = abc_11867_new_n1364
* NET 5669 = subckt_1041_nmx2_x1.q
* NET 5670 = mos6502_op[1]
* NET 5671 = abc_11867_auto_rtlil_cc_2608_muxgate_11700
* NET 5680 = abc_11867_new_n435
* NET 5682 = abc_11867_new_n1396
* NET 5683 = subckt_1662_sff1_x4.sff_s
* NET 5685 = subckt_1662_sff1_x4.y
* NET 5687 = subckt_1662_sff1_x4.sff_m
* NET 5688 = subckt_1662_sff1_x4.u
* NET 5690 = subckt_1662_sff1_x4.ckr
* NET 5691 = subckt_1662_sff1_x4.nckr
* NET 5693 = abc_11867_new_n1230
* NET 5695 = abc_11867_new_n1251
* NET 5701 = abc_11867_new_n1296
* NET 5704 = abc_11867_auto_rtlil_cc_2608_muxgate_11682
* NET 5706 = abc_11867_new_n1254
* NET 5710 = abc_11867_new_n1190
* NET 5712 = abc_11867_new_n1261
* NET 5718 = abc_11867_new_n558
* NET 5720 = abc_11867_new_n468
* NET 5724 = abc_11867_new_n1276
* NET 5728 = abc_11867_new_n1244
* NET 5730 = abc_11867_new_n469
* NET 5732 = abc_11867_new_n745
* NET 5737 = abc_11867_new_n721
* NET 5740 = abc_11867_new_n439
* NET 5817 = abc_11867_new_n1017
* NET 5823 = abc_11867_new_n1524
* NET 5825 = abc_11867_new_n1523
* NET 5828 = abc_11867_new_n912
* NET 5830 = abc_11867_new_n898
* NET 5831 = spare_buffer_11.q
* NET 5832 = spare_buffer_10.q
* NET 5833 = do[6]
* NET 5835 = abc_11867_auto_rtlil_cc_2608_muxgate_11812
* NET 5837 = abc_11867_new_n996
* NET 5838 = abc_11867_new_n945
* NET 5842 = abc_11867_new_n1377
* NET 5846 = abc_11867_flatten_mos6502_0_adj_bcd_0_0
* NET 5854 = abc_11867_new_n1354
* NET 5858 = abc_11867_new_n1235
* NET 5862 = abc_11867_new_n1187
* NET 5863 = reset_root_bl_0
* NET 5864 = clk_root_bl_2
* NET 5865 = abc_11867_new_n1229
* NET 5866 = abc_11867_new_n1208
* NET 5867 = abc_11867_new_n804
* NET 5868 = abc_11867_new_n465
* NET 5869 = abc_11867_new_n1250
* NET 5870 = abc_11867_new_n1245
* NET 5872 = abc_11867_new_n1311
* NET 5875 = abc_11867_new_n695
* NET 5876 = abc_11867_new_n461
* NET 5878 = abc_11867_new_n443
* NET 5879 = abc_11867_new_n446
* NET 5880 = di[6]
* NET 5881 = subckt_97_nmx2_x1.q
* NET 5886 = abc_11867_new_n1541
* NET 5887 = subckt_1696_sff1_x4.sff_s
* NET 5888 = mos6502_dihold[6]
* NET 5889 = subckt_1696_sff1_x4.y
* NET 5890 = subckt_1696_sff1_x4.sff_m
* NET 5891 = subckt_1696_sff1_x4.u
* NET 5892 = subckt_1696_sff1_x4.ckr
* NET 5893 = subckt_1696_sff1_x4.nckr
* NET 5896 = abc_11867_new_n1522
* NET 5897 = abc_11867_new_n1507
* NET 5898 = mos6502_pc[1]
* NET 5900 = abc_11867_new_n910
* NET 5902 = abc_11867_new_n897
* NET 5905 = abc_11867_new_n937
* NET 5906 = mos6502_pc[8]
* NET 5907 = abc_11867_new_n586
* NET 5908 = abc_11867_new_n481
* NET 5909 = abc_11867_new_n1460
* NET 5910 = abc_11867_new_n1485
* NET 5911 = abc_11867_new_n1483
* NET 5912 = abc_11867_new_n995
* NET 5913 = abc_11867_new_n993
* NET 5916 = abc_11867_new_n432
* NET 5917 = abc_11867_new_n896
* NET 5919 = abc_11867_new_n1359
* NET 5922 = abc_11867_new_n1376
* NET 5923 = abc_11867_new_n1379
* NET 5927 = abc_11867_new_n1355
* NET 5929 = abc_11867_new_n1350
* NET 5930 = subckt_1677_sff1_x4.sff_s
* NET 5931 = subckt_1677_sff1_x4.ckr
* NET 5932 = subckt_1677_sff1_x4.y
* NET 5933 = subckt_1677_sff1_x4.sff_m
* NET 5934 = subckt_1677_sff1_x4.u
* NET 5935 = abc_11867_auto_rtlil_cc_2608_muxgate_11714
* NET 5936 = subckt_1677_sff1_x4.nckr
* NET 5937 = abc_11867_new_n1264
* NET 5938 = mos6502_adc_bcd
* NET 5939 = abc_11867_new_n1265
* NET 5940 = mos6502_state[3]
* NET 5942 = abc_11867_new_n430_hfns_1
* NET 5944 = abc_11867_new_n1274
* NET 5946 = subckt_1669_sff1_x4.sff_s
* NET 5947 = subckt_1669_sff1_x4.y
* NET 5948 = subckt_1669_sff1_x4.sff_m
* NET 5949 = subckt_1669_sff1_x4.u
* NET 5950 = subckt_1669_sff1_x4.ckr
* NET 5951 = subckt_1669_sff1_x4.nckr
* NET 5952 = subckt_1678_sff1_x4.sff_s
* NET 5954 = subckt_1678_sff1_x4.y
* NET 5955 = subckt_1678_sff1_x4.sff_m
* NET 5957 = subckt_1678_sff1_x4.u
* NET 5958 = subckt_1678_sff1_x4.ckr
* NET 5960 = subckt_1678_sff1_x4.nckr
* NET 5961 = reset_root_0
* NET 5967 = abc_11867_new_n1246
* NET 5968 = abc_11867_new_n460
* NET 5971 = abc_11867_new_n1255
* NET 6008 = subckt_1737_sff1_x4.y
* NET 6010 = subckt_1737_sff1_x4.sff_m
* NET 6011 = subckt_1737_sff1_x4.ckr
* NET 6015 = abc_11867_new_n1360
* NET 6019 = abc_11867_new_n1352
* NET 6022 = subckt_1679_sff1_x4.y
* NET 6024 = subckt_1679_sff1_x4.sff_m
* NET 6025 = subckt_1679_sff1_x4.ckr
* NET 6027 = subckt_1668_sff1_x4.y
* NET 6029 = subckt_1668_sff1_x4.sff_m
* NET 6030 = subckt_1668_sff1_x4.ckr
* NET 6038 = subckt_1737_sff1_x4.sff_s
* NET 6040 = subckt_1737_sff1_x4.u
* NET 6041 = subckt_1737_sff1_x4.nckr
* NET 6043 = abc_11867_auto_rtlil_cc_2608_muxgate_11822
* NET 6050 = abc_11867_new_n1528
* NET 6051 = abc_11867_new_n1525
* NET 6055 = abc_11867_new_n1508
* NET 6062 = abc_11867_new_n946
* NET 6067 = spare_buffer_9.q
* NET 6070 = abc_11867_new_n1387
* NET 6071 = abc_11867_new_n1388
* NET 6076 = mos6502_alu_out[0]
* NET 6080 = mos6502_abh[0]
* NET 6083 = abc_11867_new_n1536
* NET 6084 = abc_11867_new_n1530
* NET 6085 = abc_11867_auto_rtlil_cc_2608_muxgate_11824
* NET 6087 = abc_11867_new_n1537
* NET 6089 = abc_11867_new_n618
* NET 6090 = abc_11867_new_n886
* NET 6095 = abc_11867_new_n1380
* NET 6096 = abc_11867_new_n1381
* NET 6102 = abc_11867_new_n1356
* NET 6103 = abc_11867_new_n1361
* NET 6112 = abc_11867_new_n1353
* NET 6125 = subckt_1679_sff1_x4.sff_s
* NET 6127 = mos6502_adc_sbc
* NET 6128 = abc_11867_auto_rtlil_cc_2608_muxgate_11718
* NET 6130 = subckt_1679_sff1_x4.nckr
* NET 6131 = subckt_1679_sff1_x4.u
* NET 6132 = abc_11867_new_n1268
* NET 6133 = abc_11867_new_n1267
* NET 6137 = abc_11867_new_n1266
* NET 6138 = abc_11867_new_n1263
* NET 6141 = mos6502_clc
* NET 6142 = abc_11867_new_n325
* NET 6143 = mos6502_shift
* NET 6144 = subckt_1668_sff1_x4.sff_s
* NET 6145 = mos6502_clv
* NET 6149 = subckt_1668_sff1_x4.u
* NET 6150 = subckt_1668_sff1_x4.nckr
* NET 6152 = clk_root_0
* NET 6154 = abc_11867_new_n1227
* NET 6156 = abc_11867_new_n1222
* NET 6157 = abc_11867_new_n1226
* NET 6158 = abc_11867_new_n1220
* NET 6161 = abc_11867_new_n1223
* NET 6166 = abc_11867_new_n1218
* NET 6172 = abc_11867_new_n540
* NET 6176 = abc_11867_new_n1243
* NET 6177 = abc_11867_new_n1312
* NET 6178 = abc_11867_new_n1308
* NET 6185 = abc_11867_new_n754
* NET 6188 = abc_11867_new_n696
* NET 6189 = abc_11867_new_n753
* NET 6191 = abc_11867_new_n755
* NET 6260 = abc_11867_new_n1543
* NET 6261 = abc_11867_new_n1545
* NET 6262 = abc_11867_new_n1527
* NET 6265 = abc_11867_new_n1534
* NET 6266 = abc_11867_new_n1533
* NET 6267 = mos6502_pc[6]
* NET 6270 = abc_11867_new_n415
* NET 6271 = abc_11867_new_n414
* NET 6273 = mos6502_pc[5]
* NET 6274 = abc_11867_new_n1521
* NET 6278 = abc_11867_new_n1511
* NET 6279 = abc_11867_new_n1505
* NET 6284 = abc_11867_new_n889
* NET 6285 = abc_11867_new_n842
* NET 6286 = abc_11867_new_n844
* NET 6288 = abc_11867_new_n911
* NET 6292 = mos6502_alu_out[7]
* NET 6293 = abc_11867_new_n428_hfns_2
* NET 6294 = abc_11867_new_n1473
* NET 6295 = abc_11867_new_n1516
* NET 6297 = abc_11867_new_n1515
* NET 6298 = abc_11867_new_n1514
* NET 6300 = abc_11867_new_n940
* NET 6301 = abc_11867_new_n939
* NET 6302 = abc_11867_new_n938
* NET 6304 = abc_11867_new_n359
* NET 6307 = abc_11867_new_n1552
* NET 6308 = abc_11867_new_n1551
* NET 6309 = abc_11867_new_n1553
* NET 6311 = abc_11867_new_n490_hfns_1
* NET 6312 = abc_11867_new_n432_hfns_2
* NET 6314 = subckt_1711_sff1_x4.sff_s
* NET 6316 = subckt_1711_sff1_x4.y
* NET 6317 = subckt_1711_sff1_x4.sff_m
* NET 6319 = abc_11867_auto_rtlil_cc_2608_muxgate_11772
* NET 6321 = subckt_1711_sff1_x4.u
* NET 6322 = subckt_1711_sff1_x4.ckr
* NET 6323 = subckt_1711_sff1_x4.nckr
* NET 6325 = abc_11867_new_n1383
* NET 6329 = abc_11867_new_n1390
* NET 6332 = abc_11867_new_n1389
* NET 6334 = abc_11867_new_n1385
* NET 6335 = abc_11867_new_n1384
* NET 6340 = abc_11867_new_n1386
* NET 6341 = mos6502_c
* NET 6344 = mos6502_n
* NET 6347 = abc_11867_new_n1372
* NET 6349 = mos6502_alu_out[3]
* NET 6353 = abc_11867_new_n1373
* NET 6358 = abc_11867_new_n326
* NET 6359 = abc_11867_new_n582
* NET 6362 = abc_11867_new_n1371
* NET 6363 = abc_11867_new_n433
* NET 6364 = subckt_1048_nmx2_x1.q
* NET 6366 = subckt_1657_sff1_x4.sff_s
* NET 6367 = subckt_1657_sff1_x4.y
* NET 6369 = subckt_1657_sff1_x4.sff_m
* NET 6371 = subckt_1657_sff1_x4.u
* NET 6372 = subckt_1657_sff1_x4.ckr
* NET 6373 = subckt_1657_sff1_x4.nckr
* NET 6374 = abc_11867_auto_rtlil_cc_2608_muxgate_11696
* NET 6375 = mos6502_bit_ins
* NET 6378 = abc_11867_new_n1217
* NET 6381 = abc_11867_new_n327
* NET 6383 = abc_11867_new_n1181_hfns_1
* NET 6384 = subckt_950_nmx2_x1.q
* NET 6386 = abc_11867_auto_rtlil_cc_2608_muxgate_11716
* NET 6388 = subckt_1663_sff1_x4.sff_s
* NET 6390 = subckt_1663_sff1_x4.sff_m
* NET 6391 = subckt_1663_sff1_x4.y
* NET 6393 = subckt_1663_sff1_x4.u
* NET 6394 = subckt_1663_sff1_x4.nckr
* NET 6395 = subckt_1663_sff1_x4.ckr
* NET 6396 = abc_11867_new_n546
* NET 6398 = mos6502_sec
* NET 6399 = abc_11867_new_n1192
* NET 6400 = abc_11867_new_n1195
* NET 6401 = abc_11867_auto_rtlil_cc_2608_muxgate_11684
* NET 6403 = abc_11867_new_n1228
* NET 6404 = abc_11867_new_n1260
* NET 6407 = abc_11867_new_n1238
* NET 6409 = abc_11867_new_n1249
* NET 6410 = abc_11867_new_n1248
* NET 6412 = abc_11867_new_n1295
* NET 6415 = abc_11867_new_n1304
* NET 6417 = abc_11867_new_n1290
* NET 6418 = abc_11867_new_n1303
* NET 6421 = abc_11867_new_n535
* NET 6466 = do[5]
* NET 6469 = abc_11867_new_n1608
* NET 6472 = abc_11867_new_n1535
* NET 6473 = abc_11867_new_n1526
* NET 6477 = abc_11867_new_n1556
* NET 6478 = abc_11867_new_n1544
* NET 6480 = abc_11867_new_n1479
* NET 6481 = abc_11867_new_n1542
* NET 6484 = mos6502_pc[7]
* NET 6485 = di[5]
* NET 6488 = subckt_93_nmx2_x1.q
* NET 6489 = mos6502_pc[3]
* NET 6490 = subckt_1735_sff1_x4.sff_s
* NET 6492 = subckt_1735_sff1_x4.y
* NET 6494 = subckt_1735_sff1_x4.sff_m
* NET 6495 = abc_11867_auto_rtlil_cc_2608_muxgate_11818
* NET 6497 = subckt_1735_sff1_x4.u
* NET 6498 = subckt_1735_sff1_x4.ckr
* NET 6499 = subckt_1735_sff1_x4.nckr
* NET 6500 = abc_11867_new_n1517
* NET 6502 = abc_11867_new_n1503
* NET 6503 = abc_11867_new_n1502
* NET 6504 = abc_11867_new_n1495
* NET 6506 = mos6502_pc[2]
* NET 6508 = subckt_1734_sff1_x4.sff_s
* NET 6509 = subckt_1734_sff1_x4.y
* NET 6510 = subckt_1734_sff1_x4.sff_m
* NET 6513 = abc_11867_auto_rtlil_cc_2608_muxgate_11816
* NET 6514 = subckt_1734_sff1_x4.ckr
* NET 6515 = subckt_1734_sff1_x4.u
* NET 6516 = subckt_1734_sff1_x4.nckr
* NET 6517 = abc_11867_new_n1726
* NET 6520 = mos6502_alu_out[6]
* NET 6524 = abc_11867_new_n343
* NET 6530 = abc_11867_new_n1009
* NET 6532 = abc_11867_new_n411
* NET 6535 = abc_11867_new_n1555
* NET 6536 = abc_11867_new_n1554
* NET 6540 = abc_11867_new_n1550
* NET 6541 = mos6502_alu_out[4]
* NET 6543 = abc_11867_new_n485_hfns_0
* NET 6544 = abc_11867_new_n428_hfns_4
* NET 6549 = mos6502_alu_out[1]
* NET 6553 = abc_11867_new_n1864
* NET 6554 = abc_11867_new_n1040
* NET 6558 = subckt_1712_sff1_x4.sff_s
* NET 6559 = subckt_1712_sff1_x4.y
* NET 6560 = subckt_1712_sff1_x4.sff_m
* NET 6563 = abc_11867_auto_rtlil_cc_2608_muxgate_11774
* NET 6564 = subckt_1712_sff1_x4.u
* NET 6565 = subckt_1712_sff1_x4.ckr
* NET 6566 = subckt_1712_sff1_x4.nckr
* NET 6567 = mos6502_z
* NET 6576 = mos6502_d
* NET 6577 = subckt_1710_sff1_x4.sff_s
* NET 6579 = subckt_1710_sff1_x4.y
* NET 6581 = abc_11867_auto_rtlil_cc_2608_muxgate_11770
* NET 6583 = subckt_1710_sff1_x4.sff_m
* NET 6584 = subckt_1710_sff1_x4.ckr
* NET 6585 = subckt_1710_sff1_x4.u
* NET 6586 = abc_11867_new_n332
* NET 6587 = subckt_1710_sff1_x4.nckr
* NET 6588 = abc_11867_new_n705
* NET 6590 = abc_11867_new_n706
* NET 6594 = abc_11867_new_n345
* NET 6597 = abc_11867_new_n707
* NET 6598 = abc_11867_new_n708
* NET 6600 = abc_11867_auto_rtlil_cc_2608_muxgate_11672
* NET 6602 = mos6502_cond_code[0]
* NET 6607 = abc_11867_new_n1370
* NET 6609 = abc_11867_new_n478_hfns_1
* NET 6614 = abc_11867_new_n1210
* NET 6615 = abc_11867_new_n1214
* NET 6617 = abc_11867_auto_rtlil_cc_2608_muxgate_11694
* NET 6618 = mos6502_plp
* NET 6620 = subckt_1660_sff1_x4.sff_s
* NET 6622 = subckt_1660_sff1_x4.y
* NET 6624 = subckt_1660_sff1_x4.sff_m
* NET 6625 = subckt_1660_sff1_x4.ckr
* NET 6626 = subckt_1660_sff1_x4.u
* NET 6627 = abc_11867_new_n1182
* NET 6628 = subckt_1660_sff1_x4.nckr
* NET 6629 = abc_11867_new_n1183
* NET 6630 = abc_11867_auto_rtlil_cc_2608_muxgate_11678
* NET 6632 = abc_11867_new_n538
* NET 6636 = abc_11867_new_n674
* NET 6639 = abc_11867_new_n676
* NET 6642 = abc_11867_new_n1232
* NET 6647 = abc_11867_new_n545
* NET 6648 = abc_11867_new_n1282
* NET 6652 = abc_11867_new_n675
* NET 6654 = abc_11867_new_n1188
* NET 6655 = abc_11867_new_n1294
* NET 6658 = abc_11867_new_n1247
* NET 6663 = abc_11867_new_n464
* NET 6667 = abc_11867_new_n751
* NET 6668 = abc_11867_new_n1310
* NET 6670 = abc_11867_new_n1309
* NET 6672 = abc_11867_new_n534_hfns_1
* NET 6754 = subckt_1743_sff1_x4.sff_s
* NET 6755 = subckt_1743_sff1_x4.y
* NET 6758 = subckt_1743_sff1_x4.sff_m
* NET 6759 = subckt_1743_sff1_x4.u
* NET 6760 = subckt_1743_sff1_x4.ckr
* NET 6761 = subckt_1743_sff1_x4.nckr
* NET 6763 = abc_11867_new_n1002
* NET 6768 = subckt_1736_sff1_x4.sff_s
* NET 6770 = subckt_1736_sff1_x4.y
* NET 6772 = subckt_1736_sff1_x4.sff_m
* NET 6773 = subckt_1736_sff1_x4.u
* NET 6774 = subckt_1736_sff1_x4.ckr
* NET 6775 = mos6502_pc[4]
* NET 6776 = subckt_1736_sff1_x4.nckr
* NET 6778 = abc_11867_new_n1518
* NET 6779 = abc_11867_new_n1513
* NET 6780 = abc_11867_auto_rtlil_cc_2608_muxgate_11820
* NET 6781 = abc_11867_new_n1519
* NET 6783 = abc_11867_new_n1510
* NET 6784 = abc_11867_new_n1501
* NET 6785 = abc_11867_new_n1492
* NET 6786 = abc_11867_new_n1509
* NET 6788 = abc_11867_new_n1748
* NET 6792 = mos6502_alu_out[5]
* NET 6793 = abc_11867_new_n342
* NET 6794 = abc_11867_new_n1085
* NET 6796 = abc_11867_new_n428_hfns_3
* NET 6797 = abc_11867_new_n485_hfns_1
* NET 6798 = abc_11867_new_n1793
* NET 6801 = mos6502_alu_out[2]
* NET 6802 = abc_11867_new_n490_hfns_0
* NET 6803 = abc_11867_new_n410
* NET 6804 = di[4]
* NET 6808 = subckt_89_nmx2_x1.q
* NET 6809 = abc_11867_new_n1770
* NET 6812 = abc_11867_new_n1818
* NET 6816 = abc_11867_new_n1070
* NET 6820 = abc_11867_new_n1073
* NET 6821 = abc_11867_new_n339
* NET 6823 = mos6502_v
* NET 6824 = subckt_1708_sff1_x4.sff_s
* NET 6826 = subckt_1708_sff1_x4.y
* NET 6827 = subckt_1708_sff1_x4.sff_m
* NET 6829 = abc_11867_auto_rtlil_cc_2608_muxgate_11764
* NET 6830 = subckt_1708_sff1_x4.u
* NET 6832 = subckt_1708_sff1_x4.nckr
* NET 6833 = subckt_1708_sff1_x4.ckr
* NET 6834 = abc_11867_new_n1843
* NET 6835 = abc_11867_new_n1672
* NET 6838 = mos6502_cond_code[2]
* NET 6840 = subckt_1659_sff1_x4.sff_s
* NET 6841 = subckt_1659_sff1_x4.y
* NET 6843 = abc_11867_auto_rtlil_cc_2608_muxgate_11676
* NET 6845 = subckt_1659_sff1_x4.sff_m
* NET 6846 = subckt_1659_sff1_x4.u
* NET 6847 = subckt_1659_sff1_x4.nckr
* NET 6848 = subckt_1659_sff1_x4.ckr
* NET 6850 = abc_11867_new_n424
* NET 6855 = subckt_1658_sff1_x4.sff_s
* NET 6856 = subckt_1658_sff1_x4.y
* NET 6859 = subckt_1658_sff1_x4.sff_m
* NET 6860 = subckt_1658_sff1_x4.u
* NET 6861 = subckt_1658_sff1_x4.ckr
* NET 6862 = subckt_1658_sff1_x4.nckr
* NET 6863 = abc_11867_auto_rtlil_cc_2608_muxgate_11674
* NET 6864 = mos6502_cond_code[1]
* NET 6867 = abc_11867_new_n330
* NET 6870 = mos6502_cld
* NET 6872 = subckt_1664_sff1_x4.sff_s
* NET 6873 = subckt_1664_sff1_x4.y
* NET 6876 = subckt_1664_sff1_x4.sff_m
* NET 6877 = subckt_1664_sff1_x4.u
* NET 6878 = subckt_1664_sff1_x4.nckr
* NET 6879 = subckt_1664_sff1_x4.ckr
* NET 6880 = abc_11867_new_n1197
* NET 6882 = abc_11867_auto_rtlil_cc_2608_muxgate_11686
* NET 6883 = mos6502_load_reg
* NET 6885 = subckt_1698_sff1_x4.sff_s
* NET 6886 = subckt_1698_sff1_x4.y
* NET 6889 = subckt_1698_sff1_x4.sff_m
* NET 6890 = subckt_1698_sff1_x4.u
* NET 6891 = subckt_1698_sff1_x4.nckr
* NET 6892 = subckt_1698_sff1_x4.ckr
* NET 6893 = abc_11867_new_n437
* NET 6897 = abc_11867_new_n1323
* NET 6899 = abc_11867_auto_rtlil_cc_2608_muxgate_11742
* NET 6900 = abc_11867_new_n441
* NET 6905 = abc_11867_new_n1224
* NET 6906 = abc_11867_new_n1225
* NET 6907 = abc_11867_new_n462
* NET 6909 = abc_11867_new_n1198
* NET 6912 = abc_11867_new_n743
* NET 6914 = abc_11867_new_n672
* NET 6915 = abc_11867_new_n1326
* NET 6917 = abc_11867_new_n1289
* NET 6918 = abc_11867_new_n673
* NET 6920 = abc_11867_new_n454
* NET 6921 = abc_11867_new_n534_hfns_0
* NET 6964 = subckt_1742_sff1_x4.sff_s
* NET 6965 = subckt_1742_sff1_x4.y
* NET 6967 = subckt_1742_sff1_x4.sff_m
* NET 6969 = subckt_1742_sff1_x4.ckr
* NET 6970 = subckt_1742_sff1_x4.u
* NET 6971 = subckt_1742_sff1_x4.nckr
* NET 6972 = abc_11867_new_n407
* NET 6974 = mos6502_dihold[5]
* NET 6976 = subckt_1695_sff1_x4.sff_s
* NET 6977 = subckt_1695_sff1_x4.y
* NET 6979 = subckt_1695_sff1_x4.sff_m
* NET 6981 = subckt_1695_sff1_x4.u
* NET 6982 = subckt_1695_sff1_x4.ckr
* NET 6983 = subckt_1695_sff1_x4.nckr
* NET 6985 = abc_11867_new_n406
* NET 6987 = di[3]
* NET 6988 = abc_11867_new_n408
* NET 6991 = subckt_85_nmx2_x1.q
* NET 6992 = mos6502_dihold[3]
* NET 6994 = subckt_1693_sff1_x4.sff_s
* NET 6995 = subckt_1693_sff1_x4.y
* NET 6998 = subckt_1693_sff1_x4.sff_m
* NET 6999 = subckt_1693_sff1_x4.ckr
* NET 7000 = subckt_1693_sff1_x4.u
* NET 7001 = subckt_1693_sff1_x4.nckr
* NET 7002 = abc_11867_new_n1639
* NET 7006 = abc_11867_new_n1627
* NET 7007 = abc_11867_new_n1626
* NET 7011 = abc_11867_new_n1638
* NET 7012 = abc_11867_new_n1092
* NET 7017 = abc_11867_new_n1628
* NET 7020 = abc_11867_new_n340
* NET 7025 = abc_11867_new_n1078
* NET 7026 = abc_11867_new_n478_hfns_0
* NET 7029 = abc_11867_new_n338
* NET 7033 = abc_11867_new_n1591
* NET 7034 = abc_11867_new_n1589
* NET 7038 = abc_11867_new_n1588
* NET 7041 = abc_11867_new_n432_hfns_1
* NET 7043 = abc_11867_new_n1590
* NET 7048 = abc_11867_new_n1064
* NET 7051 = abc_11867_new_n428_hfns_1
* NET 7053 = abc_11867_new_n1071
* NET 7056 = abc_11867_new_n337
* NET 7058 = abc_11867_new_n971
* NET 7059 = abc_11867_new_n334
* NET 7061 = abc_11867_new_n412
* NET 7062 = abc_11867_new_n1050
* NET 7065 = subckt_81_nmx2_x1.q
* NET 7068 = abc_11867_new_n986
* NET 7073 = abc_11867_new_n420
* NET 7076 = abc_11867_new_n377
* NET 7079 = subckt_1707_sff1_x4.sff_s
* NET 7080 = subckt_1707_sff1_x4.y
* NET 7082 = subckt_1707_sff1_x4.sff_m
* NET 7084 = subckt_1707_sff1_x4.u
* NET 7085 = subckt_1707_sff1_x4.ckr
* NET 7086 = subckt_1707_sff1_x4.nckr
* NET 7095 = mos6502_sed
* NET 7097 = subckt_1665_sff1_x4.sff_s
* NET 7098 = subckt_1665_sff1_x4.y
* NET 7101 = subckt_1665_sff1_x4.sff_m
* NET 7102 = subckt_1665_sff1_x4.ckr
* NET 7103 = subckt_1665_sff1_x4.u
* NET 7104 = abc_11867_new_n1202
* NET 7105 = subckt_1665_sff1_x4.nckr
* NET 7106 = abc_11867_new_n1200
* NET 7108 = abc_11867_auto_rtlil_cc_2608_muxgate_11688
* NET 7110 = abc_11867_new_n1189
* NET 7112 = abc_11867_new_n393
* NET 7114 = abc_11867_new_n1194
* NET 7119 = abc_11867_new_n392
* NET 7121 = abc_11867_new_n1216
* NET 7126 = abc_11867_new_n1234
* NET 7130 = abc_11867_new_n447
* NET 7135 = abc_11867_new_n1242
* NET 7137 = abc_11867_new_n467
* NET 7140 = abc_11867_new_n1270
* NET 7147 = abc_11867_new_n1212
* NET 7148 = abc_11867_new_n1293
* NET 7149 = abc_11867_new_n440
* NET 7151 = abc_11867_new_n627
* NET 7158 = abc_11867_new_n1241
* NET 7241 = abc_11867_auto_rtlil_cc_2608_muxgate_11832
* NET 7247 = mos6502_pc[10]
* NET 7250 = abc_11867_new_n1640
* NET 7252 = abc_11867_new_n1587
* NET 7257 = abc_11867_new_n1072
* NET 7263 = abc_11867_new_n399
* NET 7264 = abc_11867_new_n398
* NET 7270 = abc_11867_new_n378
* NET 7271 = abc_11867_auto_rtlil_cc_2608_muxgate_11762
* NET 7272 = mos6502_irhold[7]
* NET 7280 = abc_11867_new_n416
* NET 7283 = abc_11867_new_n544
* NET 7296 = abc_11867_new_n1233
* NET 7297 = abc_11867_new_n1335
* NET 7299 = abc_11867_new_n752
* NET 7300 = abc_11867_new_n1334
* NET 7301 = abc_11867_new_n1199
* NET 7302 = abc_11867_new_n1302
* NET 7304 = abc_11867_new_n1324
* NET 7305 = abc_11867_new_n541
* NET 7309 = abc_11867_new_n1582
* NET 7310 = abc_11867_new_n1584
* NET 7311 = abc_11867_new_n1573
* NET 7313 = abc_11867_new_n1583
* NET 7314 = rdy_hfns_0
* NET 7316 = abc_11867_new_n1580
* NET 7318 = abc_11867_new_n1558
* NET 7319 = abc_11867_new_n1616
* NET 7321 = abc_11867_new_n1629
* NET 7322 = abc_11867_new_n1625
* NET 7323 = abc_11867_new_n1611
* NET 7325 = abc_11867_new_n1615
* NET 7327 = abc_11867_new_n1614
* NET 7328 = abc_11867_new_n1613
* NET 7329 = abc_11867_new_n1612
* NET 7330 = abc_11867_new_n1599
* NET 7332 = abc_11867_new_n1603
* NET 7333 = abc_11867_new_n1576
* NET 7334 = abc_11867_new_n1575
* NET 7336 = abc_11867_new_n1577
* NET 7338 = abc_11867_new_n1601
* NET 7339 = abc_11867_new_n1600
* NET 7340 = abc_11867_new_n1602
* NET 7342 = abc_11867_new_n1057
* NET 7343 = abc_11867_new_n619_hfns_0
* NET 7344 = subckt_1694_sff1_x4.sff_s
* NET 7345 = mos6502_dihold[4]
* NET 7346 = subckt_1694_sff1_x4.y
* NET 7347 = subckt_1694_sff1_x4.sff_m
* NET 7348 = subckt_1694_sff1_x4.u
* NET 7349 = mos6502_dimux[4]
* NET 7350 = subckt_1694_sff1_x4.ckr
* NET 7351 = subckt_1694_sff1_x4.nckr
* NET 7352 = abc_11867_new_n432_hfns_0
* NET 7353 = abc_11867_new_n428_hfns_0
* NET 7354 = abc_11867_new_n478_hfns_2
* NET 7356 = abc_11867_new_n485_hfns_2
* NET 7357 = abc_11867_new_n1056
* NET 7358 = abc_11867_new_n1058
* NET 7359 = abc_11867_new_n1059
* NET 7361 = abc_11867_new_n436
* NET 7367 = abc_11867_new_n1049
* NET 7368 = abc_11867_new_n1051
* NET 7369 = abc_11867_new_n1052
* NET 7378 = subckt_1704_sff1_x4.sff_s
* NET 7379 = mos6502_irhold[4]
* NET 7380 = subckt_1704_sff1_x4.y
* NET 7381 = subckt_1704_sff1_x4.sff_m
* NET 7382 = subckt_1704_sff1_x4.nckr
* NET 7383 = subckt_1704_sff1_x4.u
* NET 7384 = abc_11867_auto_rtlil_cc_2608_muxgate_11756
* NET 7385 = subckt_1704_sff1_x4.ckr
* NET 7388 = subckt_1703_sff1_x4.sff_s
* NET 7389 = subckt_1703_sff1_x4.ckr
* NET 7390 = subckt_1703_sff1_x4.nckr
* NET 7391 = subckt_1703_sff1_x4.y
* NET 7392 = subckt_1703_sff1_x4.sff_m
* NET 7393 = subckt_1703_sff1_x4.u
* NET 7398 = abc_11867_new_n543
* NET 7399 = abc_11867_new_n1327
* NET 7400 = abc_11867_new_n1325
* NET 7403 = abc_11867_new_n542
* NET 7405 = abc_11867_new_n1280
* NET 7406 = do[4]
* NET 7408 = abc_11867_new_n438
* NET 7458 = abc_11867_new_n1630
* NET 7459 = abc_11867_new_n1087
* NET 7460 = abc_11867_new_n1074
* NET 7464 = abc_11867_new_n1060
* NET 7467 = subckt_1692_sff1_x4.y
* NET 7468 = subckt_1692_sff1_x4.sff_m
* NET 7470 = subckt_1692_sff1_x4.ckr
* NET 7471 = abc_11867_new_n1053
* NET 7474 = subckt_1706_sff1_x4.y
* NET 7475 = subckt_1706_sff1_x4.sff_m
* NET 7477 = subckt_1706_sff1_x4.ckr
* NET 7478 = abc_11867_new_n451
* NET 7480 = abc_11867_new_n1570
* NET 7481 = abc_11867_new_n1561
* NET 7484 = abc_11867_new_n1586
* NET 7485 = abc_11867_auto_rtlil_cc_2608_muxgate_11834
* NET 7486 = abc_11867_new_n1596
* NET 7489 = abc_11867_new_n1617
* NET 7490 = abc_11867_new_n1595
* NET 7492 = abc_11867_auto_rtlil_cc_2608_muxgate_11830
* NET 7497 = abc_11867_new_n1605
* NET 7500 = rdy_hfns_3
* NET 7503 = abc_11867_new_n1568
* NET 7508 = abc_11867_new_n1641
* NET 7512 = abc_11867_new_n1637
* NET 7513 = mos6502_pc[11]
* NET 7514 = abc_11867_new_n1624
* NET 7517 = abc_11867_new_n1592
* NET 7518 = abc_11867_new_n1593
* NET 7520 = abc_11867_new_n1578
* NET 7523 = abc_11867_new_n1574
* NET 7525 = abc_11867_new_n1086
* NET 7528 = mos6502_dimux[6]
* NET 7529 = abc_11867_new_n1084
* NET 7536 = abc_11867_new_n978
* NET 7541 = abc_11867_new_n1564
* NET 7542 = abc_11867_new_n1565
* NET 7543 = abc_11867_new_n1563
* NET 7547 = abc_11867_new_n994
* NET 7548 = abc_11867_new_n472
* NET 7549 = mos6502_dimux[7]
* NET 7550 = abc_11867_new_n507
* NET 7554 = abc_11867_new_n402
* NET 7557 = subckt_1692_sff1_x4.sff_s
* NET 7558 = mos6502_dihold[2]
* NET 7559 = abc_11867_new_n601
* NET 7561 = subckt_1692_sff1_x4.nckr
* NET 7562 = subckt_1692_sff1_x4.u
* NET 7563 = subckt_77_nmx2_x1.q
* NET 7566 = abc_11867_new_n1048
* NET 7570 = subckt_1706_sff1_x4.sff_s
* NET 7572 = mos6502_irhold[6]
* NET 7574 = subckt_1706_sff1_x4.nckr
* NET 7575 = abc_11867_auto_rtlil_cc_2608_muxgate_11760
* NET 7576 = subckt_1706_sff1_x4.u
* NET 7581 = abc_11867_new_n379
* NET 7585 = mos6502_dimux[5]
* NET 7591 = abc_11867_new_n400
* NET 7596 = abc_11867_new_n390
* NET 7603 = abc_11867_auto_rtlil_cc_2608_muxgate_11754
* NET 7604 = mos6502_irhold[3]
* NET 7612 = abc_11867_new_n404
* NET 7619 = abc_11867_new_n452
* NET 7622 = abc_11867_new_n1272
* NET 7627 = abc_11867_new_n1271
* NET 7630 = abc_11867_new_n444
* NET 7633 = abc_11867_new_n741
* NET 7639 = abc_11867_new_n1240
* NET 7643 = abc_11867_new_n453
* NET 7645 = abc_11867_new_n534_hfns_2
* NET 7646 = abc_11867_new_n534
* NET 7723 = abc_11867_new_n1571
* NET 7724 = abc_11867_new_n1557
* NET 7725 = abc_11867_new_n1569
* NET 7728 = abc_11867_new_n1607
* NET 7729 = abc_11867_new_n1618
* NET 7730 = abc_11867_new_n1594
* NET 7733 = abc_11867_new_n1633
* NET 7734 = abc_11867_new_n1631
* NET 7737 = abc_11867_new_n1604
* NET 7738 = abc_11867_new_n1606
* NET 7741 = abc_11867_new_n1645
* NET 7742 = abc_11867_new_n1632
* NET 7743 = abc_11867_new_n1644
* NET 7744 = abc_11867_new_n1635
* NET 7747 = abc_11867_new_n1477
* NET 7748 = abc_11867_new_n1579
* NET 7749 = abc_11867_new_n1581
* NET 7750 = abc_11867_new_n360
* NET 7752 = mos6502_pc[9]
* NET 7753 = abc_11867_new_n1642
* NET 7754 = abc_11867_new_n1643
* NET 7758 = abc_11867_new_n367
* NET 7759 = abc_11867_new_n1636
* NET 7760 = abc_11867_new_n1462
* NET 7761 = abc_11867_new_n1475
* NET 7765 = abc_11867_new_n1055
* NET 7766 = abc_11867_new_n361
* NET 7767 = abc_11867_new_n1094
* NET 7768 = abc_11867_new_n1091
* NET 7772 = abc_11867_new_n1088
* NET 7773 = abc_11867_new_n1083
* NET 7774 = abc_11867_new_n1093
* NET 7777 = mos6502_dimux[3]
* NET 7778 = abc_11867_new_n963
* NET 7779 = abc_11867_new_n964
* NET 7782 = abc_11867_new_n1080
* NET 7783 = abc_11867_new_n1077
* NET 7787 = abc_11867_new_n968_hfns_0
* NET 7788 = abc_11867_new_n480
* NET 7789 = abc_11867_new_n1079
* NET 7791 = abc_11867_new_n970
* NET 7793 = abc_11867_new_n1567
* NET 7794 = abc_11867_new_n1566
* NET 7796 = abc_11867_new_n1562
* NET 7797 = abc_11867_new_n1472
* NET 7798 = abc_11867_new_n576
* NET 7801 = abc_11867_new_n1069
* NET 7802 = abc_11867_new_n364
* NET 7803 = di[2]
* NET 7804 = abc_11867_new_n403
* NET 7806 = subckt_1690_sff1_x4.sff_s
* NET 7807 = subckt_1690_sff1_x4.y
* NET 7810 = subckt_1690_sff1_x4.sff_m
* NET 7811 = subckt_1690_sff1_x4.u
* NET 7812 = subckt_1690_sff1_x4.ckr
* NET 7813 = subckt_1690_sff1_x4.nckr
* NET 7814 = subckt_1727_sff1_x4.sff_s
* NET 7817 = subckt_1727_sff1_x4.y
* NET 7818 = subckt_1727_sff1_x4.sff_m
* NET 7820 = subckt_1727_sff1_x4.u
* NET 7821 = clk_root_bl_1
* NET 7822 = subckt_1727_sff1_x4.ckr
* NET 7823 = subckt_1727_sff1_x4.nckr
* NET 7824 = mos6502_abh[2]
* NET 7826 = subckt_1726_sff1_x4.sff_s
* NET 7827 = subckt_1726_sff1_x4.y
* NET 7829 = abc_11867_auto_rtlil_cc_2608_muxgate_11800
* NET 7831 = subckt_1726_sff1_x4.sff_m
* NET 7832 = subckt_1726_sff1_x4.ckr
* NET 7833 = subckt_1726_sff1_x4.nckr
* NET 7834 = subckt_1726_sff1_x4.u
* NET 7835 = mos6502_dihold[1]
* NET 7837 = subckt_1691_sff1_x4.sff_s
* NET 7838 = subckt_1691_sff1_x4.y
* NET 7841 = subckt_1691_sff1_x4.sff_m
* NET 7842 = subckt_1691_sff1_x4.u
* NET 7843 = subckt_1691_sff1_x4.ckr
* NET 7844 = subckt_1691_sff1_x4.nckr
* NET 7845 = mos6502_irhold[5]
* NET 7846 = subckt_1705_sff1_x4.sff_s
* NET 7848 = subckt_1705_sff1_x4.y
* NET 7849 = subckt_1705_sff1_x4.sff_m
* NET 7851 = abc_11867_auto_rtlil_cc_2608_muxgate_11758
* NET 7853 = subckt_1705_sff1_x4.u
* NET 7854 = subckt_1705_sff1_x4.ckr
* NET 7855 = subckt_1705_sff1_x4.nckr
* NET 7858 = abc_11867_new_n389
* NET 7863 = mos6502_dimux[1]
* NET 7867 = mos6502_irhold_valid
* NET 7869 = abc_11867_new_n435_hfns_3
* NET 7871 = abc_11867_new_n1181_hfns_0
* NET 7872 = abc_11867_new_n1193
* NET 7874 = abc_11867_new_n1213
* NET 7875 = abc_11867_new_n1329
* NET 7876 = abc_11867_new_n448
* NET 7877 = abc_11867_new_n742
* NET 7878 = abc_11867_new_n1328
* NET 7880 = abc_11867_new_n1180
* NET 7881 = abc_11867_new_n537
* NET 7882 = abc_11867_new_n539
* NET 7883 = abc_11867_new_n435_hfns_1
* NET 7884 = abc_11867_new_n463
* NET 7885 = abc_11867_new_n456
* NET 7887 = abc_11867_new_n455
* NET 7888 = abc_11867_new_n449
* NET 7889 = abc_11867_new_n1284
* NET 7890 = abc_11867_new_n1330
* NET 7891 = abc_11867_new_n435_hfns_0
* NET 7892 = abc_11867_new_n536
* NET 7893 = abc_11867_new_n442
* NET 7954 = mos6502_pc[13]
* NET 7955 = abc_11867_new_n365
* NET 7956 = abc_11867_new_n1623
* NET 7957 = rdy_hfns_2
* NET 7960 = abc_11867_new_n1610
* NET 7962 = abc_11867_new_n1620
* NET 7963 = abc_11867_auto_rtlil_cc_2608_muxgate_11838
* NET 7965 = abc_11867_new_n1619
* NET 7966 = abc_11867_new_n1621
* NET 7969 = subckt_1746_sff1_x4.sff_s
* NET 7970 = di[1]
* NET 7971 = subckt_1746_sff1_x4.y
* NET 7973 = subckt_1746_sff1_x4.sff_m
* NET 7975 = abc_11867_auto_rtlil_cc_2608_muxgate_11840
* NET 7976 = subckt_1746_sff1_x4.ckr
* NET 7977 = subckt_1746_sff1_x4.u
* NET 7978 = subckt_1746_sff1_x4.nckr
* NET 7979 = mos6502_pc[15]
* NET 7980 = subckt_1747_sff1_x4.sff_s
* NET 7982 = subckt_1747_sff1_x4.y
* NET 7984 = subckt_1747_sff1_x4.sff_m
* NET 7985 = abc_11867_auto_rtlil_cc_2608_muxgate_11842
* NET 7986 = subckt_1747_sff1_x4.u
* NET 7988 = subckt_1747_sff1_x4.ckr
* NET 7989 = subckt_1747_sff1_x4.nckr
* NET 7991 = subckt_1731_sff1_x4.sff_s
* NET 7992 = subckt_1731_sff1_x4.y
* NET 7995 = subckt_1731_sff1_x4.sff_m
* NET 7996 = subckt_1731_sff1_x4.u
* NET 7997 = subckt_1731_sff1_x4.ckr
* NET 7998 = subckt_1731_sff1_x4.nckr
* NET 7999 = abc_11867_auto_rtlil_cc_2608_muxgate_11810
* NET 8000 = mos6502_abh[7]
* NET 8004 = abc_11867_new_n1090
* NET 8006 = abc_11867_new_n1095
* NET 8008 = mos6502_pc[14]
* NET 8009 = abc_11867_new_n366
* NET 8010 = subckt_1730_sff1_x4.sff_s
* NET 8012 = subckt_1730_sff1_x4.y
* NET 8014 = subckt_1730_sff1_x4.sff_m
* NET 8015 = a[15]
* NET 8016 = subckt_1730_sff1_x4.u
* NET 8018 = subckt_1730_sff1_x4.ckr
* NET 8019 = subckt_1730_sff1_x4.nckr
* NET 8020 = abc_11867_auto_rtlil_cc_2608_muxgate_11808
* NET 8021 = mos6502_abh[6]
* NET 8025 = abc_11867_new_n1076
* NET 8028 = abc_11867_new_n1081
* NET 8030 = subckt_1729_sff1_x4.sff_s
* NET 8031 = subckt_1729_sff1_x4.y
* NET 8034 = subckt_1729_sff1_x4.sff_m
* NET 8035 = subckt_1729_sff1_x4.ckr
* NET 8036 = subckt_1729_sff1_x4.u
* NET 8037 = subckt_1729_sff1_x4.nckr
* NET 8038 = a[14]
* NET 8039 = abc_11867_auto_rtlil_cc_2608_muxgate_11806
* NET 8040 = mos6502_abh[5]
* NET 8045 = abc_11867_new_n954_hfns_0
* NET 8046 = abc_11867_new_n362
* NET 8047 = abc_11867_new_n968_hfns_1
* NET 8048 = abc_11867_new_n975
* NET 8051 = abc_11867_new_n395
* NET 8052 = abc_11867_new_n1063
* NET 8053 = abc_11867_new_n1065
* NET 8054 = abc_11867_new_n1066
* NET 8055 = di[0]
* NET 8058 = abc_11867_new_n396
* NET 8059 = mos6502_dihold[0]
* NET 8061 = abc_11867_new_n394
* NET 8062 = subckt_73_nmx2_x1.q
* NET 8063 = clk_root_br_0
* NET 8064 = rdy_hfns_1
* NET 8066 = a[13]
* NET 8067 = abc_11867_new_n1067
* NET 8068 = abc_11867_new_n1062
* NET 8070 = abc_11867_auto_rtlil_cc_2608_muxgate_11802
* NET 8071 = mos6502_abh[3]
* NET 8077 = subckt_1728_sff1_x4.sff_s
* NET 8078 = subckt_1728_sff1_x4.y
* NET 8079 = subckt_1728_sff1_x4.sff_m
* NET 8082 = subckt_1728_sff1_x4.u
* NET 8083 = subckt_1728_sff1_x4.ckr
* NET 8084 = subckt_1728_sff1_x4.nckr
* NET 8085 = abc_11867_auto_rtlil_cc_2608_muxgate_11804
* NET 8086 = mos6502_abh[4]
* NET 8089 = a[12]
* NET 8094 = abc_11867_new_n1443
* NET 8097 = mos6502_abh[1]
* NET 8099 = subckt_1725_sff1_x4.sff_s
* NET 8100 = subckt_1725_sff1_x4.y
* NET 8102 = abc_11867_auto_rtlil_cc_2608_muxgate_11798
* NET 8104 = subckt_1725_sff1_x4.sff_m
* NET 8105 = subckt_1725_sff1_x4.ckr
* NET 8106 = subckt_1725_sff1_x4.u
* NET 8107 = subckt_1725_sff1_x4.nckr
* NET 8109 = a[11]
* NET 8110 = subckt_1700_sff1_x4.sff_s
* NET 8111 = subckt_1700_sff1_x4.y
* NET 8113 = subckt_1700_sff1_x4.sff_m
* NET 8115 = subckt_1700_sff1_x4.u
* NET 8116 = subckt_1700_sff1_x4.ckr
* NET 8117 = subckt_1700_sff1_x4.nckr
* NET 8118 = abc_11867_auto_rtlil_cc_2608_muxgate_11748
* NET 8119 = mos6502_irhold[0]
* NET 8122 = mos6502_dimux[0]
* NET 8125 = mos6502_irhold[1]
* NET 8127 = subckt_1701_sff1_x4.sff_s
* NET 8128 = subckt_1701_sff1_x4.y
* NET 8130 = abc_11867_auto_rtlil_cc_2608_muxgate_11750
* NET 8132 = subckt_1701_sff1_x4.sff_m
* NET 8133 = subckt_1701_sff1_x4.u
* NET 8134 = subckt_1701_sff1_x4.ckr
* NET 8135 = subckt_1701_sff1_x4.nckr
* NET 8136 = a[10]
* NET 8137 = abc_11867_new_n391
* NET 8139 = mos6502_dimux[2]
* NET 8140 = abc_11867_new_n1341
* NET 8144 = vdd
* NET 8145 = abc_11867_new_n435_hfns_4
* NET 8147 = mos6502_irhold[2]
* NET 8148 = subckt_1702_sff1_x4.sff_s
* NET 8150 = subckt_1702_sff1_x4.y
* NET 8152 = subckt_1702_sff1_x4.sff_m
* NET 8153 = abc_11867_auto_rtlil_cc_2608_muxgate_11752
* NET 8154 = subckt_1702_sff1_x4.u
* NET 8156 = a[9]
* NET 8157 = subckt_1702_sff1_x4.ckr
* NET 8158 = subckt_1702_sff1_x4.nckr
* NET 8159 = mos6502_store
* NET 8161 = subckt_1683_sff1_x4.sff_s
* NET 8162 = subckt_1683_sff1_x4.y
* NET 8165 = subckt_1683_sff1_x4.sff_m
* NET 8166 = clk_root_bl_0
* NET 8167 = subckt_1683_sff1_x4.ckr
* NET 8168 = subckt_1683_sff1_x4.u
* NET 8169 = abc_11867_new_n1287
* NET 8170 = subckt_1683_sff1_x4.nckr
* NET 8171 = abc_11867_new_n1285
* NET 8172 = abc_11867_new_n1286
* NET 8173 = abc_11867_auto_rtlil_cc_2608_muxgate_11726
* NET 8175 = abc_11867_new_n1331
* NET 8176 = abc_11867_new_n1333
* NET 8179 = abc_11867_new_n1211
* NET 8180 = abc_11867_new_n1301
* NET 8182 = abc_11867_new_n1332
* NET 8184 = abc_11867_new_n435_hfns_2
* NET 8185 = vss
* NET 8186 = abc_11867_new_n450
* NET 8187 = abc_11867_new_n445
* NET 8188 = abc_11867_new_n466
Mtr_16868 8144 7336 7335 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16867 7335 7333 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16866 8144 7334 7335 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16865 7520 7335 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16864 8144 662 659 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16863 662 923 587 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16862 586 663 662 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16861 8144 923 663 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16860 587 3537 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16859 8144 676 586 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16858 659 662 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16857 8144 258 256 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16856 258 923 218 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16855 217 260 258 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16854 8144 923 260 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16853 218 3532 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16852 8144 266 217 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16851 256 258 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16850 3378 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16849 3378 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16848 8144 4293 3378 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16847 8144 6896 6893 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16846 6896 7867 6895 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16845 6894 6898 6896 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16844 8144 7867 6898 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16843 6895 7061 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16842 8144 7112 6894 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16841 6893 6896 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16840 8144 7117 7408 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16839 7117 7867 6945 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16838 6944 7120 7117 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16837 8144 7867 7120 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16836 6945 7349 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16835 8144 7379 6944 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16834 7408 7117 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16833 1583 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16832 1583 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16831 8144 5654 1583 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16830 8144 7051 1583 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16829 8144 1455 1291 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16828 1291 1710 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16827 8144 1729 1291 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16826 1293 1291 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16825 3674 3722 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16824 3718 3717 3674 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16823 8144 3971 3718 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16822 6650 7140 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16821 8144 7147 6650 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16820 6648 6650 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16819 6124 7361 5999 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16818 5999 6907 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16817 8144 6576 6124 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16816 6133 6124 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16815 7873 8179 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16814 8144 7872 7873 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16813 7874 7873 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16812 3976 4009 3977 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16811 3974 7787 3976 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16810 3975 8048 3974 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16809 8144 8045 3975 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16808 3972 3977 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16807 8144 4574 2824 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16806 2824 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16805 2824 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16804 8144 6484 2824 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16803 2822 2824 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16802 5142 5440 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16801 8144 5139 5142 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16800 5140 5142 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16799 8144 1284 62 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16798 4644 1928 63 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16797 63 1284 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16796 63 62 4644 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16795 8144 61 63 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16794 61 1928 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16793 7482 7723 7409 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16792 8144 7481 7409 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16791 7409 7480 7482 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16790 7492 7482 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16789 2445 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16788 8144 5942 2445 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16787 2894 2445 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16786 941 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16785 8144 5654 941 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16784 1352 941 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16783 4692 5406 4591 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16782 4591 6821 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16781 8144 6809 4692 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16780 4690 4692 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16779 561 562 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16778 762 764 561 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16777 8144 1364 762 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16776 4741 4738 4601 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16775 4601 4737 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16774 8144 4739 4741 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16773 4983 4741 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16772 8144 6156 5696 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16771 5696 6157 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16770 5696 6166 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16769 8144 7880 5696 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16768 5695 5696 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16767 5056 8047 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16766 5154 5907 5056 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16765 8144 6541 5154 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16764 2948 4470 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16763 8144 3033 2948 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16762 2947 2948 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16761 8144 6797 4930 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16760 4930 7026 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16759 8144 6544 4930 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16758 5907 4930 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16757 5742 7408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16756 8144 7883 5742 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16755 5740 5742 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16754 8144 3405 3178 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16753 3178 3177 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16752 3178 4276 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16751 8144 3404 3178 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16750 3872 3178 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16749 8144 4068 2008 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16748 2008 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16747 8144 2492 2008 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16746 2006 2008 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16745 8144 559 167 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16744 167 558 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16743 8144 1362 167 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16742 166 167 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16741 4446 4535 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16740 4444 4532 4531 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16739 8144 4720 4444 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16738 4532 4536 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16737 8144 5864 4536 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16736 8144 4721 4535 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16735 4534 4532 4446 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16734 4445 4536 4534 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16733 8144 4533 4445 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16732 4533 4534 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16731 4531 4536 4533 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16730 8144 4531 4720 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16729 4720 4531 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16728 8144 6802 5626 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16727 5626 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16726 8144 5624 5626 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16725 7798 5626 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16724 1588 1891 1013 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16723 1012 2698 1588 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16722 8144 1996 1012 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16721 1013 2926 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16720 8144 7398 6397 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16719 6397 6907 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16718 8144 7891 6397 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16717 6396 6397 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16716 8144 5654 2257 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16715 2257 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16714 2257 5483 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16713 8144 3857 2257 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16712 2256 2257 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16711 8144 4051 3397 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16710 3397 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16709 3397 7026 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16708 8144 5624 3397 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16707 3635 3397 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16706 2330 2344 2276 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16705 2276 2601 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16704 8144 2589 2330 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16703 2596 2330 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16702 8144 6152 5904 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16701 5832 5904 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16700 8144 5904 5832 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16699 8144 5904 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16698 8144 5904 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16697 8144 5961 5903 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16696 5831 5903 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16695 8144 5903 5831 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16694 8144 5903 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16693 8144 5903 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16692 8144 6152 2021 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16691 3834 2021 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16690 8144 2021 3834 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16689 8144 2021 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16688 8144 2021 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16687 8144 6152 2020 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16686 2019 2020 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16685 8144 2020 2019 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16684 8144 2020 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16683 8144 2020 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16682 8144 6152 1810 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16681 1809 1810 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16680 8144 1810 1809 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16679 8144 1810 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16678 8144 1810 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16677 8144 5961 1808 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16676 1807 1808 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16675 8144 1808 1807 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16674 8144 1808 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16673 8144 1808 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16672 8144 6152 1953 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16671 3708 1953 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16670 8144 1953 3708 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16669 8144 1953 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16668 8144 1953 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16667 8144 6152 1952 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16666 1951 1952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16665 8144 1952 1951 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16664 8144 1952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16663 8144 1952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16662 8144 6152 1748 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16661 1772 1748 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16660 8144 1748 1772 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16659 8144 1748 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16658 8144 1748 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16657 8144 5961 1747 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16656 1746 1747 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16655 8144 1747 1746 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16654 8144 1747 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16653 8144 1747 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16652 6002 6178 6001 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16651 6001 6668 6181 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16650 6181 6672 6002 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16649 6002 7151 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16648 8144 6658 6002 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16647 6177 6181 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16646 8144 190 189 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16645 188 189 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16644 8144 1699 188 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16643 187 188 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16642 8144 188 187 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16641 8144 2041 1873 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16640 1873 2039 3182 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16639 482 483 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16638 477 484 478 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16637 8144 676 477 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16636 484 485 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16635 8144 1951 485 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16634 8144 659 483 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16633 480 484 482 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16632 481 485 480 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16631 8144 479 481 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16630 479 480 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16629 478 485 479 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16628 8144 478 676 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16627 676 478 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16626 6931 7000 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16625 6929 6999 6994 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16624 8144 6992 6929 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16623 6999 7001 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16622 8144 8063 7001 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16621 8144 7777 7000 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16620 6998 6999 6931 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16619 6930 7001 6998 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16618 8144 6995 6930 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16617 6995 6998 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16616 6994 7001 6995 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16615 8144 6994 6992 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16614 6992 6994 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16613 1474 3969 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16612 8144 1473 1474 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16611 1003 1115 1004 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16610 1004 1114 1109 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16609 1109 1113 1004 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16608 1003 1111 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16607 8144 1110 1003 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16606 1004 1116 1003 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16605 1325 1109 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16604 7411 7490 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16603 7965 7497 7411 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16602 8144 7489 7965 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16601 2796 7549 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16600 2796 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16599 8144 4172 2796 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16598 6936 7084 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16597 6934 7085 7079 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16596 8144 7272 6934 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16595 7085 7086 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16594 8144 7821 7086 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16593 8144 7271 7084 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16592 7082 7085 6936 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16591 6935 7086 7082 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16590 8144 7080 6935 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16589 7080 7082 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16588 7079 7086 7080 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16587 8144 7079 7272 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16586 7272 7079 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16585 7781 7778 7780 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16584 7780 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16583 8144 7777 7781 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16582 8052 7781 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16581 8136 7464 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16580 8144 7765 8136 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16579 3267 3186 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16578 8144 3187 3267 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16577 1000 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16576 1158 2227 1000 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16575 999 1157 1158 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16574 8144 2698 999 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16573 2022 1158 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16572 4954 6090 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16571 4953 6089 4954 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16570 8144 6341 4953 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16569 7898 7977 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16568 7896 7976 7969 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16567 8144 8008 7896 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16566 7976 7978 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16565 8144 8063 7978 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16564 8144 7975 7977 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16563 7973 7976 7898 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16562 7897 7978 7973 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16561 8144 7971 7897 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16560 7971 7973 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16559 7969 7978 7971 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16558 8144 7969 8008 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16557 8008 7969 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16556 5504 5503 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16555 5504 5507 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16554 8144 5508 5504 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16553 8144 7880 5504 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16552 7110 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16551 7110 7892 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16550 8144 7408 7110 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16549 957 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16548 8144 7051 957 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16547 8144 1588 1437 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16546 1435 1589 1902 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16545 1436 1587 1435 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16544 1437 1892 1436 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16543 8144 1616 1439 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16542 1440 1617 1816 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16541 1441 1618 1440 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16540 1439 1615 1441 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16539 3103 3543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16538 8144 3553 3103 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16537 3102 3103 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16536 6320 6321 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16535 6315 6322 6314 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16534 8144 6344 6315 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16533 6322 6323 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16532 8144 8063 6323 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16531 8144 6319 6321 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16530 6317 6322 6320 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16529 6318 6323 6317 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16528 8144 6316 6318 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16527 6316 6317 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16526 6314 6323 6316 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16525 8144 6314 6344 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16524 6344 6314 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16523 2666 2669 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16522 2662 2670 2663 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16521 8144 6076 2662 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16520 2670 2671 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16519 8144 3708 2671 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16518 8144 2668 2669 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16517 2667 2670 2666 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16516 2665 2671 2667 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16515 8144 2664 2665 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16514 2664 2667 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16513 2663 2671 2664 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16512 8144 2663 6076 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16511 6076 2663 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16510 6053 6778 5978 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16509 5978 6051 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16508 8144 7314 6053 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16507 6050 6053 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16506 5427 5629 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16505 8144 5426 5427 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16504 5618 5427 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16503 5536 5641 5535 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16502 5535 5653 5639 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16501 5639 5642 5536 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16500 5536 5637 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16499 8144 5644 5536 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16498 6095 5639 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16497 5508 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16496 5508 6909 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16495 8144 6636 5508 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16494 8144 7130 5508 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16493 6629 7130 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16492 6629 7880 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16491 8144 6921 6629 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16490 8156 7471 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16489 8144 7566 8156 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16488 7876 8184 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16487 7876 7630 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16486 8144 7893 7876 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16485 8144 3356 3138 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16484 3138 3579 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16483 8144 3582 3138 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16482 3137 3138 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16481 1295 1729 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16480 1295 1455 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16479 8144 1710 1295 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16478 1299 5395 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16477 8144 1301 1299 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16476 1719 1299 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16475 3755 4511 3683 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16474 8144 4510 3683 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16473 3683 4512 3755 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16472 3754 3755 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16471 3331 3763 3210 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16470 8144 4510 3210 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16469 3210 4424 3331 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16468 3330 3331 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16467 5028 5504 5029 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16466 5029 6177 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16465 8144 5026 5028 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16464 5027 5028 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16463 5249 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16462 5249 8179 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16461 8144 6654 5249 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16460 8144 7130 5249 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16459 5693 6158 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16458 5693 5865 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16457 8144 6154 5693 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16456 6403 6632 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16455 6403 6906 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16454 8144 6647 6403 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16453 2467 3172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16452 2467 2238 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16451 8144 2239 2467 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16450 5499 5503 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16449 8144 7880 5499 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16448 5500 5499 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16447 6905 8184 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16446 6905 7398 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16445 8144 7881 6905 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16444 8144 4900 4670 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16443 4672 7029 4588 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16442 4588 4900 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16441 4588 4670 4672 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16440 8144 4671 4588 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16439 4671 7029 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16438 3654 4078 3653 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16437 3652 3851 3654 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16436 8144 3651 3652 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16435 3650 3653 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16434 8144 3073 3074 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16433 3074 3650 3194 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16432 3197 3194 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16431 7886 7889 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16430 8144 7885 7886 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16429 8171 7886 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16428 8144 7121 6169 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16427 6169 6652 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16426 8144 6636 6169 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16425 6378 6169 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16424 7516 7760 7418 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16423 7418 7761 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16422 8144 8008 7516 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16421 7514 7516 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16420 8144 3577 3578 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16419 4502 3575 3576 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16418 3576 3577 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16417 3576 3578 4502 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16416 8144 3574 3576 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16415 3574 3575 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16414 8144 3175 2921 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16413 7353 2921 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16412 8144 2921 7353 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16411 8144 2921 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16410 8144 2921 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16409 8144 3175 781 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16408 7051 781 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16407 8144 781 7051 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16406 8144 781 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16405 8144 781 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16404 8144 3175 3176 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16403 6293 3176 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16402 8144 3176 6293 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16401 8144 3176 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16400 8144 3176 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16399 8144 3175 2457 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16398 6796 2457 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16397 8144 2457 6796 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16396 8144 2457 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16395 8144 2457 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16394 8144 3175 3169 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16393 6544 3169 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16392 8144 3169 6544 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16391 8144 3169 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16390 8144 3169 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16389 8144 369 368 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16388 3175 368 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16387 8144 368 3175 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16386 8144 368 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16385 8144 368 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16384 8144 3844 3174 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16383 3174 4295 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16382 3172 3399 3174 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16381 3173 3170 3172 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16380 3174 3171 3173 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16379 3870 3867 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16378 8144 4292 3870 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16377 3868 3870 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16376 8144 1184 1183 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16375 3857 1183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16374 8144 1183 3857 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16373 8144 1183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16372 8144 1183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16371 8144 1184 1185 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16370 4075 1185 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16369 8144 1185 4075 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16368 8144 1185 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16367 8144 1185 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16366 8144 963 964 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16365 1184 964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16364 8144 964 1184 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16363 8144 964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16362 8144 964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16361 8144 6775 6779 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16360 8144 7500 6777 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16359 6779 6777 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16358 8144 365 160 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16357 160 553 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16356 8144 166 160 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16355 334 160 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16354 8144 7026 2197 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16353 2197 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16352 2197 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16351 8144 6080 2197 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16350 2198 2197 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16349 8144 2896 2770 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16348 2770 4067 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16347 7058 6796 2770 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16346 2769 2898 7058 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16345 2770 2894 2769 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16344 8144 2485 2487 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16343 2487 2484 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16342 8144 2947 2487 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16341 2955 2487 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16340 4686 5406 4589 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16339 4589 7029 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16338 8144 6798 4686 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16337 4685 4686 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16336 5857 5949 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16335 5855 5950 5946 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16334 8144 6375 5855 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16333 5950 5951 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16332 8144 7821 5951 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16331 8144 6374 5949 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16330 5948 5950 5857 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16329 5856 5951 5948 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16328 8144 5947 5856 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16327 5947 5948 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16326 5946 5951 5947 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16325 8144 5946 6375 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16324 6375 5946 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16323 5073 5238 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16322 5226 6629 5073 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16321 8144 5223 5226 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16320 8144 4895 4654 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16319 4663 6524 4586 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16318 4586 4895 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16317 4586 4654 4663 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16316 8144 4655 4586 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16315 4655 6524 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16314 8144 7026 1380 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16313 1380 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16312 1380 5624 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16311 8144 3857 1380 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16310 1593 1380 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16309 8144 4068 1179 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16308 1179 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16307 1179 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16306 8144 3857 1179 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16305 2252 1179 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16304 3586 3783 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16303 8144 3782 3586 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16302 3212 3774 3211 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16301 3211 3587 3342 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16300 3342 3579 3212 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16299 3212 3780 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16298 8144 4255 3212 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16297 3340 3342 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16296 208 304 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16295 206 303 298 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16294 8144 709 206 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16293 303 305 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16292 8144 1772 305 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16291 8144 710 304 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16290 302 303 208 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16289 207 305 302 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16288 8144 299 207 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16287 299 302 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16286 298 305 299 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16285 8144 298 709 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16284 709 298 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16283 5063 5193 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16282 5061 5195 5186 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16281 8144 5197 5061 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16280 5195 5194 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16279 8144 5864 5194 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16278 8144 5196 5193 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16277 5191 5195 5063 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16276 5062 5194 5191 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16275 8144 5189 5062 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16274 5189 5191 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16273 5186 5194 5189 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16272 8144 5186 5197 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16271 5197 5186 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16270 5438 6294 5439 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16269 5439 7059 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16268 8144 5437 5438 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16267 5436 5438 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16266 6015 6520 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16265 8144 6618 6015 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16264 6614 6383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16263 8144 6145 6614 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16262 4580 5037 4475 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16261 4475 4583 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16260 8144 4579 4580 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16259 4474 4580 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16258 4115 4583 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16257 4315 5041 4115 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16256 8144 4317 4315 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16255 3423 3419 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16254 8144 3264 3423 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16253 3782 3780 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16252 8144 4543 3782 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16251 2813 5401 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16250 8144 2159 2813 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16249 3122 3569 3124 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16248 3124 3123 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16247 8144 3567 3122 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16246 3121 3122 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16245 5866 7872 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16244 8144 6396 5866 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16243 5489 6383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16242 8144 5485 5489 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16241 5494 6654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16240 8144 6396 5494 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16239 5486 6383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16238 8144 5202 5486 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16237 5739 5879 5546 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16236 5546 7887 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16235 8144 5878 5739 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16234 5737 5739 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16233 3664 3871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16232 8144 3665 3664 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16231 3264 3268 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16230 8144 3192 3264 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16229 553 1150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16228 8144 6363 553 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16227 5829 5898 5827 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16226 5902 7752 5829 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16225 5829 6285 5902 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16224 5827 6286 5829 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16223 5827 6549 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16222 8144 6284 5827 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16221 1929 1924 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16220 8144 1711 1929 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16219 7830 7834 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16218 7825 7832 7826 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16217 8144 7824 7825 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16216 7832 7833 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16215 8144 8166 7833 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16214 8144 7829 7834 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16213 7831 7832 7830 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16212 7828 7833 7831 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16211 8144 7827 7828 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16210 7827 7831 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16209 7826 7833 7827 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16208 8144 7826 7824 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16207 7824 7826 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16206 5388 5387 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16205 5388 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16204 8144 7352 5388 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16203 619 955 761 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16202 618 762 619 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16201 8144 956 618 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16200 943 761 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16199 6949 7029 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16198 8054 7058 6949 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16197 8144 7048 8054 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16196 1559 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16195 1559 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16194 8144 4573 1559 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16193 5868 7884 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16192 8144 8184 5868 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16191 4288 5031 4111 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16190 4111 4583 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16189 8144 4286 4288 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16188 4287 4288 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_16187 7324 7325 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16186 8144 7323 7324 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16185 7319 7324 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16184 3140 3146 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16183 8144 4007 3140 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16182 3139 3140 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16181 7909 8016 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16180 7907 8018 8010 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16179 8144 8021 7907 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16178 8018 8019 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16177 8144 8063 8019 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_16176 8144 8020 8016 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16175 8014 8018 7909 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16174 7908 8019 8014 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16173 8144 8012 7908 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16172 8012 8014 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16171 8010 8019 8012 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16170 8144 8010 8021 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16169 8021 8010 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16168 5452 5665 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_16167 5455 8122 5451 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16166 5451 6359 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16165 8144 5450 5457 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16164 5457 5658 5454 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16163 5454 5452 5455 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16162 5455 5665 5456 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16161 5456 5453 5457 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16160 8144 6359 5450 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_16159 5449 5455 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16158 8144 495 496 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16157 495 923 452 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16156 451 453 495 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16155 8144 923 453 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16154 452 3978 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16153 8144 497 451 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16152 496 495 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16151 8144 921 920 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16150 921 923 924 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16149 922 925 921 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16148 8144 923 925 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16147 924 4012 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16146 8144 1111 922 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16145 920 921 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16144 8144 698 697 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16143 698 923 599 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16142 598 701 698 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16141 8144 923 701 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16140 599 4160 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16139 8144 703 598 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16138 697 698 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16137 8144 728 724 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16136 728 923 608 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16135 607 727 728 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16134 8144 923 727 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16133 608 4176 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16132 8144 725 607 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16131 724 728 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16130 8144 290 287 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16129 290 923 226 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16128 225 291 290 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16127 8144 923 291 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16126 226 3999 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16125 8144 512 225 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16124 287 290 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16123 5168 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16122 5168 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16121 8144 4573 5168 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16120 1368 2013 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16119 8144 3148 1368 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16118 7328 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16117 7328 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16116 8144 6797 7328 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16115 8144 6792 7328 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16114 2165 2166 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16113 8144 3229 2165 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16112 2355 2165 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16111 7253 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16110 7252 7798 7253 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16109 8144 7777 7252 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16108 8144 5628 5433 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16107 5433 5629 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16106 8144 5434 5433 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16105 5432 5433 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16104 8144 307 306 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16103 307 923 230 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16102 229 310 307 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16101 8144 923 310 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16100 230 2402 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16099 8144 529 229 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16098 306 307 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16097 8144 892 890 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16096 892 1332 893 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16095 891 894 892 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16094 8144 1332 894 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16093 893 3537 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16092 8144 1048 891 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16091 890 892 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16090 8144 1039 1038 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16089 1039 1332 979 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16088 980 1042 1039 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16087 8144 1332 1042 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16086 979 3532 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16085 8144 1043 980 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16084 1038 1039 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16083 8144 887 885 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16082 887 1332 888 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16081 886 889 887 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16080 8144 1332 889 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16079 888 3978 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16078 8144 1304 886 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16077 885 887 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16076 5110 5938 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16075 5110 6801 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16074 8144 5108 5110 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16073 8144 5606 5110 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16072 3379 5624 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16071 3379 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16070 8144 4167 3379 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16069 6191 7299 6006 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16068 6005 6188 6191 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16067 8144 6667 6005 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16066 6006 6189 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16065 2245 2941 2244 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16064 2243 2241 2245 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16063 8144 2242 2243 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16062 3656 2244 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16061 3804 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16060 3804 4167 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16059 8144 5447 3804 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16058 8144 5664 3804 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16057 8144 4173 2811 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16056 2811 4172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16055 8144 7528 2811 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16054 2809 2811 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16053 8144 3744 1836 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16052 1836 2602 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16051 1924 2141 1836 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16050 1835 3737 1924 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16049 1836 2136 1835 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16048 1893 1887 1804 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16047 1803 2698 1893 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16046 8144 6359 1803 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16045 1804 2926 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_16044 6806 6808 7061 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16043 8144 7500 6808 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_16042 6807 7345 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16041 7061 7500 6807 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16040 8144 6804 6806 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16039 2782 2941 2945 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16038 2781 2942 2782 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16037 8144 2946 2781 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_16036 3645 2945 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16035 2367 2379 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_16034 2370 3562 2286 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16033 2286 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16032 8144 2364 2288 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16031 2288 2365 2287 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16030 2287 2367 2370 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16029 2370 2379 2289 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16028 2289 2843 2288 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16027 8144 3556 2364 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_16026 2635 2370 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16025 2357 2379 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_16024 2358 2352 2282 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16023 2282 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16022 8144 2353 2284 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16021 2284 2355 2283 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16020 2283 2357 2358 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16019 2358 2379 2285 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16018 2285 2840 2284 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_16017 8144 3556 2353 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_16016 3108 2358 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16015 8144 4197 4199 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16014 8047 4199 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16013 8144 4199 8047 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16012 8144 4199 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16011 8144 4199 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16010 8144 3771 3772 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16009 4197 3772 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16008 8144 3772 4197 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16007 8144 3772 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16006 8144 3772 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16005 8144 5654 5650 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16004 5650 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16003 5650 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16002 8144 6375 5650 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_16001 5929 5650 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_16000 6426 6488 7280 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15999 8144 7500 6488 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15998 6425 6974 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15997 7280 7500 6425 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15996 8144 6485 6426 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15995 7953 8186 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15994 8188 8187 7953 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15993 8144 8184 8188 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15992 366 1150 235 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15991 235 3391 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15990 8144 3393 366 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15989 365 366 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15988 5901 5902 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15987 8144 5917 5901 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15986 5830 5901 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15985 1347 1348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15984 8144 1346 1347 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15983 4025 1347 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15982 8144 4197 4008 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15981 7787 4008 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15980 8144 4008 7787 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15979 8144 4008 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15978 8144 4008 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15977 8144 5108 5105 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15976 5121 5938 5051 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15975 5051 5108 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15974 5051 5105 5121 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15973 8144 5102 5051 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15972 5102 5938 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15971 5818 7559 5816 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15970 5816 7548 5884 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15969 5884 7550 5818 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15968 5818 6270 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15967 8144 6271 5818 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15966 5817 5884 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15965 499 1115 500 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15964 500 1114 501 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15963 501 685 500 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15962 499 497 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15961 8144 1110 499 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15960 500 498 499 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15959 1738 501 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15958 6810 6835 6811 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15957 6811 7061 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15956 8144 7053 6810 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15955 6809 6810 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15954 2632 2631 2634 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15953 2634 2836 2633 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15952 2633 3744 2634 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15951 2632 2636 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15950 8144 3112 2632 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15949 2634 2630 2632 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15948 2830 2633 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15947 8144 2133 1286 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15946 1284 2132 1285 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15945 1285 2133 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15944 1285 1286 1284 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15943 8144 1283 1285 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15942 1283 2132 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15941 8144 4951 4711 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15940 7343 4711 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15939 8144 4711 7343 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15938 8144 4711 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15937 8144 4711 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15936 8144 4951 4952 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15935 5574 4952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15934 8144 4952 5574 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15933 8144 4952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15932 8144 4952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15931 8144 4525 4526 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15930 4951 4526 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15929 8144 4526 4951 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15928 8144 4526 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15927 8144 4526 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15926 8144 6403 5964 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15925 5964 6156 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15924 8144 6166 5964 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15923 5865 5964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15922 7377 7398 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15921 8144 7891 7377 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15920 7283 7377 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15919 2606 3320 2607 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15918 2607 2809 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15917 8144 3315 2606 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15916 2605 2606 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15915 3555 3748 3554 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15914 3554 3552 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15913 8144 3553 3555 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15912 3740 3555 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15911 3810 3809 3688 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15910 3688 3812 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15909 8144 7314 3810 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15908 4737 3810 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15907 6436 6524 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15906 7767 7058 6436 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15905 8144 7012 7767 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15904 5376 7559 5375 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15903 5375 7548 5374 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15902 5374 7550 5376 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15901 5376 5373 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15900 8144 5551 5376 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15899 5372 5374 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15898 1367 1570 1366 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15897 1366 1571 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15896 8144 1364 1367 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15895 1365 1367 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15894 8144 2262 237 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15893 237 5940 576 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15892 3742 3740 3681 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15891 3681 3743 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15890 8144 4141 3742 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15889 4157 3742 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15888 1755 2179 1754 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15887 1754 2178 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15886 8144 1962 1755 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15885 2170 1755 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15884 3289 4492 3200 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15883 3200 3720 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15882 8144 3286 3289 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15881 3287 3289 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15880 211 318 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15879 209 317 312 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15878 8144 725 209 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15877 317 319 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15876 8144 1772 319 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15875 8144 724 318 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15874 316 317 211 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15873 210 319 316 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15872 8144 313 210 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15871 313 316 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15870 312 319 313 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15869 8144 312 725 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15868 725 312 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15867 5020 5022 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15866 5016 5023 5017 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15865 8144 5015 5016 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15864 5023 5024 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15863 8144 5864 5024 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15862 8144 5027 5022 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15861 5021 5023 5020 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15860 5019 5024 5021 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15859 8144 5018 5019 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15858 5018 5021 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15857 5017 5024 5018 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15856 8144 5017 5015 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15855 5015 5017 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15854 6462 6639 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15853 6630 6629 6462 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15852 8144 6627 6630 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15851 4598 4955 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15850 7361 4730 4598 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15849 8144 4731 7361 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15848 8144 2718 1394 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15847 1394 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15846 1394 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15845 8144 5648 1394 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15844 1616 1394 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15843 8144 3641 3643 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15842 3643 3642 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15841 3643 4299 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15840 8144 4287 3643 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15839 3660 3643 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15838 8144 5148 560 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15837 560 2203 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15836 560 1372 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15835 8144 1157 560 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15834 558 560 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15833 202 254 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15832 200 253 248 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15831 8144 266 200 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15830 253 255 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15829 8144 1951 255 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15828 8144 256 254 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15827 250 253 202 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15826 201 255 250 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15825 8144 249 201 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15824 249 250 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15823 248 255 249 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15822 8144 248 266 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15821 266 248 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15820 8144 7314 7308 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15819 7307 7308 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15818 8144 7513 7307 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15817 7484 7307 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15816 8144 7307 7484 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15815 7360 7788 7261 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15814 7261 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15813 8144 7824 7360 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15812 7358 7360 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15811 2201 2202 2412 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15810 2200 2198 2201 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15809 8144 2199 2200 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15808 8144 3603 2763 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15807 2764 2887 3009 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15806 2765 2888 2764 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15805 2763 3606 2765 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15804 2140 2141 2139 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15803 2139 2612 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15802 8144 2136 2140 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15801 2138 2140 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15800 7365 7562 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15799 7363 7470 7557 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15798 8144 7558 7363 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15797 7470 7561 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15796 8144 7821 7561 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15795 8144 8139 7562 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15794 7468 7470 7365 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15793 7364 7561 7468 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15792 8144 7467 7364 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15791 7467 7468 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15790 7557 7561 7467 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15789 8144 7557 7558 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15788 7558 7557 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15787 4885 6261 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15786 8144 8064 4885 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15785 6881 7110 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15784 6882 7106 6881 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15783 8144 6880 6882 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15782 1490 4137 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15781 8144 1315 1490 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15780 7374 7576 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15779 7372 7477 7570 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15778 8144 7572 7372 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15777 7477 7574 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15776 8144 8166 7574 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15775 8144 7575 7576 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15774 7475 7477 7374 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15773 7373 7574 7475 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15772 8144 7474 7373 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15771 7474 7475 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15770 7570 7574 7474 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15769 8144 7570 7572 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15768 7572 7570 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15767 4401 4483 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15766 4399 4484 4480 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15765 8144 7954 4399 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15764 4484 4485 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15763 8144 8063 4485 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15762 8144 7963 4483 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15761 4482 4484 4401 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15760 4400 4485 4482 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15759 8144 4481 4400 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15758 4481 4482 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15757 4480 4485 4481 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15756 8144 4480 7954 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15755 7954 4480 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15754 8182 8188 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15753 8182 8180 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15752 8144 8179 8182 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15751 7890 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15750 7890 7892 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15749 8144 7884 7890 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15748 1154 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15747 8144 2718 1154 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15746 1364 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15745 8144 4067 1364 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15744 3151 3150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15743 8144 6363 3151 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15742 3361 3151 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15741 4104 7029 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15740 4171 5406 4104 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15739 8144 6798 4171 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15738 3290 3720 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15737 8144 4492 3290 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15736 3717 3290 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15735 6450 6585 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15734 6448 6584 6577 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15733 8144 6576 6448 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15732 6584 6587 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15731 8144 7821 6587 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15730 8144 6581 6585 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15729 6583 6584 6450 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15728 6449 6587 6583 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15727 8144 6579 6449 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15726 6579 6583 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15725 6577 6587 6579 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15724 8144 6577 6576 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15723 6576 6577 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15722 8144 4571 4460 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15721 4571 7871 4462 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15720 4463 4464 4571 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15719 8144 7871 4464 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15718 4462 5030 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15717 8144 4461 4463 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15716 4460 4571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15715 6382 6384 6386 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15714 8144 6383 6384 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15713 6385 7622 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15712 6386 6383 6385 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15711 8144 6381 6382 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15710 2390 2408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15709 8144 4433 2390 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15708 8144 7729 7732 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15707 7732 7738 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15706 8144 7730 7732 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15705 7962 7732 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15704 7014 7012 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15703 8144 7343 7014 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15702 7011 7014 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15701 8144 7759 7756 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15700 7755 7756 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15699 8144 7753 7755 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15698 7754 7755 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15697 8144 7755 7754 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15696 3607 3802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15695 8144 4032 3607 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15694 3606 3607 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15693 8144 2849 2847 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15692 2849 3327 2742 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15691 2741 2851 2849 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15690 8144 3327 2851 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15689 2742 3348 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15688 8144 3315 2741 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15687 2847 2849 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15686 7240 7310 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15685 7241 7313 7240 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15684 8144 7311 7241 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15683 7404 7405 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15682 8144 7478 7404 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15681 7304 7404 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15680 1849 1964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15679 1966 1965 1849 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15678 8144 4429 1966 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15677 8144 2256 1872 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15676 1872 2258 2034 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15675 2039 2034 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15674 8144 2964 2967 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15673 2966 2967 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15672 8144 2968 2966 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15671 3662 2966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15670 8144 2966 3662 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15669 8144 3635 3638 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15668 3638 3636 3637 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15667 4070 3637 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15666 2890 2421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15665 2890 2424 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15664 8144 2430 2890 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15663 8144 4203 2890 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15662 7499 7747 7412 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15661 7412 7802 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15660 8144 7737 7499 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15659 7497 7499 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15658 4424 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15657 4424 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15656 8144 4574 4424 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15655 8144 5898 4424 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15654 8144 6658 5874 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15653 5874 7151 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15652 5872 6672 5874 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15651 5873 6668 5872 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15650 5874 6178 5873 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15649 6363 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15648 6363 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15647 8144 5942 6363 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15646 8144 7137 5545 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15645 5545 5876 5731 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15644 5730 5731 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15643 1416 1477 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15642 4927 1476 1416 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15641 8144 3148 4927 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15640 8144 1559 1556 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15639 1556 1796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15638 1556 1806 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15637 8144 1891 1556 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15636 1558 1556 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15635 8144 5169 1984 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15634 1984 4517 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15633 1984 2227 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15632 8144 4518 1984 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15631 1985 1984 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15630 8144 3109 3106 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15629 3313 3108 3110 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15628 3110 3109 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15627 3110 3106 3313 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15626 8144 3107 3110 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15625 3107 3108 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15624 6280 6278 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15623 6495 6783 6280 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15622 8144 6279 6495 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15621 3970 4648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15620 8144 3972 3970 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15619 3969 3970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15618 4442 4705 4521 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15617 4441 8047 4442 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15616 4440 8048 4441 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15615 8144 8045 4440 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15614 4439 4521 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15613 5135 5420 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15612 8144 5132 5135 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15611 5133 5135 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15610 7922 8062 8058 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15609 8144 8064 8062 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15608 7923 8059 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15607 8058 8064 7923 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15606 8144 8055 7922 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15605 8144 2492 622 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15604 622 1799 768 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15603 1800 768 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15602 2784 2962 2963 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15601 2785 3865 2784 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15600 8144 3258 2785 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15599 2961 2963 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15598 2432 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15597 8144 4068 2432 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15596 2682 2432 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15595 4519 4942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15594 8144 4945 4519 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15593 4438 4519 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15592 6303 6301 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15591 8144 6302 6303 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15590 6300 6303 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15589 1998 1999 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15588 8144 1996 1998 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15587 2424 1998 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15586 2691 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15585 8144 4167 2691 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15584 3370 2691 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15583 8144 4310 4217 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15582 4217 7354 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15581 8144 6293 4217 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15580 6089 4217 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15579 8144 3872 3873 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15578 3873 3876 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15577 8144 4479 3873 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15576 3871 3873 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15575 8144 4489 4487 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15574 4403 4651 4404 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15573 4404 4489 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15572 4404 4487 4403 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15571 8144 4488 4404 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15570 4488 4651 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15569 8144 7026 3634 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15568 3634 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15567 8144 7353 3634 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15566 3842 3634 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15565 387 2262 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15564 8144 5940 387 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15563 386 387 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15562 6800 6835 6799 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15561 6799 6988 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15560 8144 7048 6800 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15559 6798 6800 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15558 1294 1293 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15557 1298 1292 1294 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15556 8144 1954 1298 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15555 2312 2500 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15554 2310 2499 2494 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15553 8144 2492 2310 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15552 2499 2501 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15551 8144 3834 2501 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15550 8144 3661 2500 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15549 2496 2499 2312 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15548 2311 2501 2496 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15547 8144 2495 2311 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15546 2495 2496 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15545 2494 2501 2495 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15544 8144 2494 2492 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15543 2492 2494 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15542 5959 6149 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15541 5953 6030 6144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15540 8144 6145 5953 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15539 6030 6150 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15538 8144 7821 6150 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15537 8144 6617 6149 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15536 6029 6030 5959 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15535 5956 6150 6029 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15534 8144 6027 5956 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15533 6027 6029 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15532 6144 6150 6027 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15531 8144 6144 6145 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15530 6145 6144 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15529 8144 5188 3616 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15528 7314 3616 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15527 8144 3616 7314 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15526 8144 3616 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15525 8144 3616 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15524 8144 5188 3808 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15523 8064 3808 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15522 8144 3808 8064 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15521 8144 3808 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15520 8144 3808 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15519 8144 5188 5172 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15518 7957 5172 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15517 8144 5172 7957 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15516 8144 5172 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15515 8144 5172 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15514 8144 5188 5173 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15513 7500 5173 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15512 8144 5173 7500 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15511 8144 5173 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15510 8144 5173 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15509 8144 4079 4080 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15508 5188 4080 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15507 8144 4080 5188 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15506 8144 4080 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15505 8144 4080 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15504 8144 4068 1824 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15503 1824 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15502 1824 4167 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15501 8144 7353 1824 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15500 1825 1824 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15499 8144 1825 1826 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15498 1826 1827 2036 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15497 6464 6918 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15496 6667 6663 6464 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15495 8144 7149 6667 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15494 1821 4518 1374 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_15493 1373 2698 1821 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_15492 8144 1372 1373 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_15491 1374 2926 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_15490 3581 3780 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15489 8144 5197 3581 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15488 214 330 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15487 212 332 325 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15486 8144 535 212 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15485 332 333 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15484 8144 3834 333 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15483 8144 549 330 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15482 329 332 214 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15481 213 333 329 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15480 8144 327 213 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15479 327 329 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15478 325 333 327 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15477 8144 325 535 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15476 535 325 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15475 7534 7778 7428 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15474 7428 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15473 8144 7585 7534 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15472 7783 7534 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15471 8144 4293 1600 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15470 1600 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15469 1600 5483 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15468 8144 3857 1600 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15467 1898 1600 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15466 2864 2866 2759 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15465 2759 2877 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15464 8144 2863 2864 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15463 3575 2864 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15462 4453 4546 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15461 4451 4547 4542 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15460 8144 4543 4451 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15459 4547 4549 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15458 8144 5864 4549 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15457 8144 5213 4546 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15456 4545 4547 4453 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15455 4452 4549 4545 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15454 8144 4544 4452 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15453 4544 4545 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15452 4542 4549 4544 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15451 8144 4542 4543 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15450 4543 4542 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15449 5144 5143 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15448 5144 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15447 8144 7352 5144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15446 6019 6359 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15445 8144 6363 6019 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15444 7104 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15443 8144 7095 7104 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15442 6880 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15441 8144 6870 6880 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15440 3162 3787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15439 8144 3787 3160 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15438 3159 5453 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15437 8144 3159 3162 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15436 3162 3160 3161 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15435 3161 5453 3162 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15434 3158 3161 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15433 8144 3161 3158 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15432 4276 5867 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15431 8144 4790 4276 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15430 7935 8106 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15429 7933 8105 8099 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15428 8144 8097 7933 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15427 8105 8107 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15426 8144 8166 8107 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15425 8144 8102 8106 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15424 8104 8105 7935 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15423 7934 8107 8104 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15422 8144 8100 7934 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15421 8100 8104 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15420 8099 8107 8100 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15419 8144 8099 8097 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15418 8097 8099 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15417 6480 5434 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15416 6480 5628 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15415 8144 5629 6480 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15414 6400 7872 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15413 8144 6652 6400 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15412 8144 741 740 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15411 741 903 612 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15410 613 744 741 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15409 8144 903 744 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15408 612 4176 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15407 8144 739 613 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15406 740 741 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15405 8144 4179 4176 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15404 4179 4178 4087 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15403 4086 4181 4179 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15402 8144 4178 4181 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15401 4087 4925 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15400 8144 8139 4086 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15399 4176 4179 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15398 4786 7887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15397 8144 7130 4786 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15396 8144 3857 3699 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15395 3699 3844 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15394 3847 4575 3699 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15393 3698 7788 3847 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15392 3699 3842 3698 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15391 4010 4517 4011 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15390 8144 4009 4011 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15389 4011 4518 4010 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15388 4192 4010 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15387 1927 2152 1837 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15386 8144 2616 1837 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15385 1837 2608 1927 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15384 1925 1927 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15383 3992 4511 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15382 8144 4512 3992 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15381 3991 3992 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15380 1762 1760 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15379 3134 1761 1762 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15378 8144 1962 3134 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15377 3146 8122 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15376 3146 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15375 8144 4172 3146 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15374 8144 3744 2758 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15373 2758 3139 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15372 2875 3130 2758 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15371 2757 3737 2875 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15370 2758 2860 2757 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15369 5819 6524 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15368 6481 6294 5819 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15367 8144 5886 6481 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15366 5405 5414 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15365 5588 5616 5405 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15364 8144 7957 5588 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15363 7452 7877 7451 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15362 7451 7876 7623 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15361 7623 7627 7452 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15360 7452 7883 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15359 8144 7884 7452 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15358 7622 7623 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15357 5858 7126 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15356 8144 6154 5858 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15355 8144 1334 1330 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15354 1334 1332 1333 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15353 1331 1336 1334 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15352 8144 1332 1336 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15351 1333 4012 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15350 8144 1335 1331 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15349 1330 1334 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15348 8144 1077 1074 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15347 1077 1332 988 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15346 987 1078 1077 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15345 8144 1332 1078 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15344 988 4160 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15343 8144 1317 987 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15342 1074 1077 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15341 4548 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15340 4548 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15339 8144 7026 4548 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15338 5434 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15337 5434 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15336 8144 6543 5434 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15335 1887 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15334 1887 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15333 8144 7026 1887 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15332 6920 7643 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15331 8144 7869 6920 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15330 4298 7026 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15329 4298 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15328 8144 4068 4298 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15327 8144 4067 4298 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15326 4473 7887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15325 4473 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15324 8144 4790 4473 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15323 8144 5740 4473 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15322 6286 4517 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15321 8144 4518 6286 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15320 8144 7957 7961 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15319 7959 7961 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15318 8144 8008 7959 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15317 7956 7959 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15316 8144 7959 7956 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15315 3819 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15314 3819 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15313 8144 5447 3819 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15312 8144 4260 3819 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15311 2160 5401 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15310 8144 2159 2160 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15309 2619 2160 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15308 2658 2877 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15307 8144 2866 2658 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15306 2659 2658 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15305 8144 7340 7337 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15304 7337 7338 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15303 8144 7339 7337 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15302 7332 7337 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15301 8144 7749 7315 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15300 7315 7725 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15299 8144 7724 7315 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15298 7313 7315 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15297 8144 1323 1506 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15296 1323 1332 1321 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15295 1322 1324 1323 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15294 8144 1332 1324 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15293 1321 4176 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15292 8144 1499 1322 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15291 1506 1323 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15290 8144 918 915 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15289 918 1332 917 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15288 916 919 918 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15287 8144 1332 919 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15286 917 3999 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15285 8144 1088 916 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15284 915 918 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15283 8144 1094 1091 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15282 1094 1332 993 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15281 992 1096 1094 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15280 8144 1332 1096 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15279 993 2402 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15278 8144 1758 992 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15277 1091 1094 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15276 8144 897 1069 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15275 897 939 895 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15274 896 898 897 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15273 8144 939 898 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15272 895 3537 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15271 8144 1063 896 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15270 1069 897 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15269 8144 274 272 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15268 274 939 224 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15267 223 277 274 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15266 8144 939 277 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15265 224 3532 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15264 8144 273 223 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15263 272 274 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15262 5169 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15261 5169 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15260 8144 4574 5169 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15259 8144 1593 1438 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15258 1438 1597 1594 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15257 1892 1594 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15256 2821 3757 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_15255 2817 2813 2736 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15254 2736 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15253 8144 2815 2739 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15252 2739 2816 2737 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15251 2737 2821 2817 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15250 2817 3757 2738 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15249 2738 3303 2739 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15248 8144 3556 2815 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_15247 3095 2817 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15246 2623 3757 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_15245 2626 2619 2622 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15244 2622 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15243 8144 2620 2627 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15242 2627 2621 2624 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15241 2624 2623 2626 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15240 2626 3757 2625 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15239 2625 3307 2627 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15238 8144 3556 2620 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_15237 3098 2626 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15236 8144 6359 5645 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15235 5645 5908 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15234 8144 6363 5645 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15233 5644 5645 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15232 8144 502 691 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15231 502 939 455 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15230 454 456 502 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15229 8144 939 456 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15228 455 3978 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15227 8144 685 454 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15226 691 502 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15225 8144 937 935 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15224 937 939 936 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15223 938 940 937 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15222 8144 939 940 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15221 936 4012 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15220 8144 1113 938 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15219 935 937 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15218 1796 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15217 1796 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15216 8144 4572 1796 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15215 6189 6893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15214 6189 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15213 8144 7893 6189 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15212 8144 7883 6189 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15211 5041 6396 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15210 5041 5875 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15209 8144 6636 5041 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15208 8144 6921 5041 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15207 5273 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15206 5273 6652 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15205 8144 6172 5273 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15204 8144 6921 5273 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15203 8144 4529 4524 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15202 4524 4707 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15201 4524 4548 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15200 8144 4527 4524 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15199 7761 4524 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15198 4767 5501 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15197 8144 4766 4767 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15196 4765 4767 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15195 5001 5701 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15194 8144 7880 5001 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15193 5002 5001 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15192 1125 1132 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15191 8144 8064 1125 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15190 1123 1125 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15189 7713 7802 7800 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15188 7714 8047 7713 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15187 7712 8048 7714 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15186 8144 8045 7712 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_15185 7801 7800 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15184 8144 3744 3572 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15183 3572 3571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15182 3570 3569 3572 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15181 3568 3737 3570 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15180 3572 3567 3568 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15179 6290 6775 6291 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15178 8144 6295 6291 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15177 6291 6480 6290 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15176 6500 6290 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15175 4555 6383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15174 8144 4556 4555 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15173 5212 4555 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15172 8144 370 183 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15171 4310 183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15170 8144 183 4310 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15169 8144 183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15168 8144 183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15167 8144 370 371 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15166 1565 371 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15165 8144 371 1565 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15164 8144 371 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15163 8144 371 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15162 8144 185 182 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15161 370 182 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15160 8144 182 370 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15159 8144 182 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15158 8144 182 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15157 8144 1968 1763 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15156 8045 1763 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15155 8144 1763 8045 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15154 8144 1763 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15153 8144 1763 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15152 8144 1968 1969 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15151 4429 1969 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15150 8144 1969 4429 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15149 8144 1969 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15148 8144 1969 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15147 8144 1776 1764 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15146 1968 1764 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15145 8144 1764 1968 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15144 8144 1764 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15143 8144 1764 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15142 2911 4167 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15141 8144 5654 2911 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15140 3371 2911 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15139 1326 1325 1328 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15138 1328 1327 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15137 8144 1962 1326 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15136 3997 1326 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15135 6268 6267 6269 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15134 8144 6266 6269 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15133 6269 6480 6268 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15132 6472 6268 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15131 4237 6867 4110 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15130 4110 4236 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15129 8144 7867 4237 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15128 4738 4237 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15127 2302 2894 2301 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15126 2301 2898 2426 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15125 2426 6796 2302 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15124 2302 4067 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15123 8144 2896 2302 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15122 2677 2426 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15121 7585 7280 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15120 7528 7073 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15119 6649 7884 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15118 8144 8184 6649 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15117 6663 6649 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15116 8144 4575 2725 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15115 2725 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15114 2725 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15113 8144 5483 2725 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15112 2950 2725 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15111 8144 4540 1363 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15110 1363 1996 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15109 8144 1986 1363 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15108 1362 1363 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15107 8144 359 357 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15106 357 1150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15105 8144 4251 357 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15104 354 357 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15103 1912 6469 1831 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15102 8144 1909 1831 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15101 1831 7728 1912 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15100 1910 1912 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15099 8144 3744 2629 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15098 2629 2836 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15097 3109 3112 2629 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15096 2628 3737 3109 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15095 2629 3108 2628 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15094 205 284 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15093 203 285 278 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15092 8144 512 203 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15091 285 286 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15090 8144 1951 286 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15089 8144 287 284 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15088 282 285 205 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15087 204 286 282 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15086 8144 280 204 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15085 280 282 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15084 278 286 280 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15083 8144 278 512 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15082 512 278 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15081 4057 4059 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15080 4053 4060 4054 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15079 8144 4461 4053 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15078 4060 4062 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15077 8144 5864 4062 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15076 8144 4460 4059 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15075 4058 4060 4057 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15074 4056 4062 4058 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15073 8144 4055 4056 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15072 4055 4058 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15071 4054 4062 4055 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15070 8144 4054 4461 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15069 4461 4054 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15068 8144 4672 4500 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15067 4414 5109 4415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15066 4415 4672 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15065 4415 4500 4414 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15064 8144 4501 4415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15063 4501 5109 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_15062 8144 6609 960 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15061 960 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15060 960 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15059 8144 3857 960 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15058 1168 960 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15057 7349 7061 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15056 8144 5483 4064 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15055 4064 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15054 4064 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15053 8144 4075 4064 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15052 4790 4064 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15051 3770 5406 3685 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15050 3685 4939 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15049 8144 6553 3770 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15048 3768 3770 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15047 2598 3287 2597 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15046 2597 2596 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15045 8144 2594 2598 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15044 2595 2598 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_15043 490 492 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15042 487 493 486 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15041 8144 497 487 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15040 493 494 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15039 8144 1951 494 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15038 8144 496 492 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15037 491 493 490 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15036 488 494 491 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15035 8144 489 488 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15034 489 491 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15033 486 494 489 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15032 8144 486 497 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15031 497 486 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15030 7840 7842 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15029 7836 7843 7837 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15028 8144 7835 7836 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15027 7843 7844 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15026 8144 8166 7844 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15025 8144 7863 7842 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15024 7841 7843 7840 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15023 7839 7844 7841 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15022 8144 7838 7839 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15021 7838 7841 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15020 7837 7844 7838 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15019 8144 7837 7835 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15018 7835 7837 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15017 1978 4184 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15016 8144 1966 1978 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_15015 8144 4295 4113 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15014 4113 4997 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15013 4292 4790 4113 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15012 4112 5732 4292 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15011 4113 6912 4112 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_15010 7852 7853 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15009 7847 7854 7846 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15008 8144 7845 7847 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15007 7854 7855 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15006 8144 8166 7855 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_15005 8144 7851 7853 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15004 7849 7854 7852 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15003 7850 7855 7849 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15002 8144 7848 7850 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15001 7848 7849 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_15000 7846 7855 7848 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14999 8144 7846 7845 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14998 7845 7846 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14997 6083 6472 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14996 8144 6473 6083 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14995 2678 2677 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14994 8144 6076 2678 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14993 8144 2492 7548 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14992 8144 1799 364 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14991 7548 364 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14990 1962 1355 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14989 1962 1357 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14988 8144 1558 1962 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14987 8144 3319 3316 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14986 3319 3748 3206 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14985 3207 3321 3319 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14984 8144 3748 3321 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14983 3206 3348 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14982 8144 3315 3207 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14981 3316 3319 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14980 473 474 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14979 468 475 469 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14978 8144 3077 468 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14977 475 476 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14976 8144 3708 476 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14975 8144 1910 474 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14974 472 475 473 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14973 471 476 472 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14972 8144 470 471 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14971 470 472 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14970 469 476 470 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14969 8144 469 3077 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14968 3077 469 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14967 7040 7048 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14966 8144 7343 7040 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14965 7038 7040 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14964 8144 8003 7999 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14963 8003 8094 7906 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14962 7905 8005 8003 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14961 8144 8094 8005 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14960 7906 8015 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14959 8144 8000 7905 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14958 7999 8003 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14957 8144 8023 8020 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14956 8023 8094 7911 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14955 7910 8027 8023 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14954 8144 8094 8027 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14953 7911 8038 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14952 8144 8021 7910 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14951 8020 8023 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14950 8144 8042 8039 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14949 8042 8094 7916 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14948 7915 8044 8042 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14947 8144 8094 8044 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14946 7916 8066 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14945 8144 8040 7915 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14944 8039 8042 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14943 8144 8087 8085 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14942 8087 8094 7930 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14941 7929 8091 8087 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14940 8144 8094 8091 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14939 7930 8089 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14938 8144 8086 7929 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14937 8085 8087 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14936 8144 8074 8070 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14935 8074 8094 7925 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14934 7924 8075 8074 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14933 8144 8094 8075 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14932 7925 8109 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14931 8144 8071 7924 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14930 8070 8074 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14929 8144 7569 7829 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14928 7569 8094 7438 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14927 7437 7571 7569 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14926 8144 8094 7571 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14925 7438 8136 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14924 8144 7824 7437 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14923 7829 7569 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14922 3063 3711 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14921 8144 1047 3063 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14920 8144 4714 4701 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14919 8144 7314 4622 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14918 4701 4622 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14917 8144 1799 562 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14916 8144 2492 563 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14915 562 563 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14914 8144 2477 2026 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14913 2024 2026 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14912 8144 2022 2024 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14911 2238 2024 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14910 8144 2024 2238 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14909 2888 2205 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14908 2888 2207 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14907 8144 2206 2888 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14906 2142 2803 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14905 8144 3553 2142 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14904 2141 2142 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14903 4512 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14902 4512 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14901 8144 5648 4512 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14900 8144 6489 4512 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14899 2319 3752 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14898 8144 2318 2319 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14897 8144 6786 6787 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14896 6787 6784 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14895 8144 6785 6787 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14894 6783 6787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14893 8144 8093 8102 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14892 8093 8094 7932 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14891 7931 8096 8093 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14890 8144 8094 8096 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14889 7932 8156 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14888 8144 8097 7931 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14887 8102 8093 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14886 5701 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14885 5701 8179 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14884 8144 7872 5701 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14883 8144 7130 5701 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14882 8144 1154 954 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14881 954 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14880 954 5147 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14879 8144 1543 954 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14878 1358 954 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14877 8144 4572 4031 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14876 4031 7354 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14875 4031 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14874 8144 6143 4031 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14873 4234 4031 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14872 8144 3997 3998 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14871 3996 3998 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14870 8144 4690 3996 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14869 3995 3996 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14868 8144 3996 3995 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14867 8144 6478 6474 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14866 6474 6477 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14865 6474 6472 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14864 8144 6473 6474 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14863 7724 6474 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14862 5826 7029 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14861 6055 6294 5826 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14860 8144 5897 6055 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14859 5115 5114 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14858 8144 7056 5115 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14857 5113 5115 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14856 8144 2262 186 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14855 184 186 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14854 8144 5940 184 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14853 185 184 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14852 8144 184 185 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14851 8144 7892 7894 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14850 7894 7893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14849 8144 7891 7894 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14848 8180 7894 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14847 1759 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14846 8144 1758 1759 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14845 2178 1759 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14844 1320 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14843 8144 1499 1320 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14842 1964 1320 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14841 8144 4498 4153 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14840 4152 4149 4102 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14839 4102 4498 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14838 4102 4153 4152 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14837 8144 4150 4102 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14836 4150 4149 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14835 4132 4133 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14834 8144 4129 4132 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14833 4130 4132 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14832 3403 4075 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14831 8144 4734 3403 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14830 3399 3403 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14829 2692 4306 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14828 2913 4302 2692 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14827 8144 3371 2913 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14826 5402 5406 5403 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14825 5403 7020 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14824 8144 6788 5402 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14823 5401 5402 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14822 8144 4402 1749 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14821 4489 6793 1751 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14820 1751 4402 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14819 1751 1749 4489 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14818 8144 1750 1751 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14817 1750 6793 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14816 8144 7403 6913 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14815 6913 7881 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14814 8144 7891 6913 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14813 6918 6913 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14812 8144 3863 3864 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14811 3864 4476 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14810 8144 4299 3864 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14809 3860 3864 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14808 3196 3425 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14807 3190 3424 3421 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14806 8144 5940 3190 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14805 3424 3426 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14804 8144 3834 3426 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14803 8144 3423 3425 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14802 3271 3424 3196 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14801 3195 3426 3271 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14800 8144 3270 3195 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14799 3270 3271 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14798 3421 3426 3270 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14797 8144 3421 5940 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14796 5940 3421 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14795 8144 7957 5548 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14794 5549 5548 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14793 8144 7752 5549 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14792 7481 5549 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14791 8144 5549 7481 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14790 4757 6412 4603 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14789 4603 5002 4757 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14788 8144 4756 4603 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14787 7355 7788 7258 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14786 7258 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14785 8144 8086 7355 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14784 7257 7355 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14783 8144 2246 2248 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14782 2248 2247 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14781 8144 3172 2248 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14780 2958 2248 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14779 8144 6609 1175 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14778 1175 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14777 1175 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14776 8144 3857 1175 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14775 1173 1175 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14774 8144 7887 4783 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14773 4783 7130 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14772 8144 7149 4783 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14771 4782 4783 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14770 8144 344 337 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14769 337 352 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14768 337 551 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14767 8144 349 337 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14766 5641 337 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14765 8144 3340 2760 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14764 2760 3009 2867 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14763 2866 2867 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14762 5072 5222 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14761 5070 5221 5216 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14760 8144 5485 5070 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14759 5221 5224 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14758 8144 5864 5224 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14757 8144 5490 5222 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14756 5219 5221 5072 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14755 5071 5224 5219 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14754 8144 5217 5071 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14753 5217 5219 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14752 5216 5224 5217 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14751 8144 5216 5485 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14750 5485 5216 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14749 8144 5447 1829 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14748 1829 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14747 1829 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14746 8144 4075 1829 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14745 1904 1829 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14744 118 120 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14743 114 121 115 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14742 8144 514 114 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14741 121 122 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14740 8144 1951 122 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14739 8144 292 120 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14738 119 121 118 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14737 117 122 119 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14736 8144 116 117 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14735 116 119 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14734 115 122 116 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14733 8144 115 514 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14732 514 115 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14731 5462 5464 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14730 5458 5465 5459 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14729 8144 5670 5458 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14728 5465 5466 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14727 8144 7821 5466 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14726 8144 5671 5464 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14725 5463 5465 5462 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14724 5461 5466 5463 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14723 8144 5460 5461 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14722 5460 5463 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14721 5459 5466 5460 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14720 8144 5459 5670 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14719 5670 5459 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14718 3670 3707 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14717 3668 3710 3701 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14716 8144 3956 3668 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14715 3710 3709 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14714 8144 3708 3709 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14713 8144 3955 3707 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14712 3705 3710 3670 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14711 3669 3709 3705 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14710 8144 3703 3669 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14709 3703 3705 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14708 3701 3709 3703 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14707 8144 3701 3956 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14706 3956 3701 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14705 8140 4737 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14704 8144 4739 8140 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14703 6399 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14702 8144 6398 6399 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14701 5710 6654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14700 8144 6652 5710 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14699 3667 3877 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14698 8144 4318 3667 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14697 7740 7741 7699 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14696 8144 7744 7699 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14695 7699 7743 7740 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14694 7985 7740 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14693 8144 4770 4033 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14692 8144 6143 4034 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14691 4033 4034 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14690 3229 3348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14689 8144 3315 3229 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14688 7338 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14687 7338 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14686 8144 6543 7338 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14685 8144 6541 7338 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14684 1356 1353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14683 1356 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14682 8144 5654 1356 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14681 6899 7297 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14680 8144 6897 6899 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14679 5862 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14678 8144 6141 5862 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14677 5223 6383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14676 8144 5003 5223 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14675 8144 527 528 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14674 527 903 458 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14673 457 459 527 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14672 8144 903 459 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14671 458 3999 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14670 8144 517 457 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14669 528 527 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14668 6359 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14667 6359 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14666 8144 6543 6359 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14665 7478 8186 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14664 8144 8184 7478 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14663 4479 6191 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14662 8144 4790 4479 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14661 1822 2032 1899 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14660 1823 1821 1822 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14659 8144 2249 1823 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14658 6285 5147 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14657 8144 5148 6285 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14656 2144 5395 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14655 8144 1301 2144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14654 2298 2400 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14653 2296 2399 2393 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14652 8144 6080 2296 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14651 2399 2401 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14650 8144 3708 2401 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14649 8144 2398 2400 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14648 2397 2399 2298 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14647 2297 2401 2397 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14646 8144 2394 2297 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14645 2394 2397 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14644 2393 2401 2394 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14643 8144 2393 6080 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14642 6080 2393 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14641 7490 7725 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14640 7490 7518 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14639 8144 7749 7490 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14638 8144 7724 7490 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14637 7320 7747 7246 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14636 7246 7766 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14635 8144 7748 7320 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14634 7316 7320 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14633 8144 4002 3999 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14632 4002 4178 4000 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14631 4001 4004 4002 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14630 8144 4178 4004 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14629 4000 4698 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14628 8144 7863 4001 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14627 3999 4002 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14626 8144 144 141 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14625 144 903 142 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14624 143 145 144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14623 8144 903 145 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14622 142 2402 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14621 8144 530 143 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14620 141 144 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14619 4420 7559 4419 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14618 4419 7548 4504 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14617 4504 7550 4420 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14616 4420 4507 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14615 8144 4701 4420 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14614 4418 4504 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14613 4527 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14612 4527 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14611 8144 4051 4527 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14610 8144 7558 7554 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14609 8144 7957 7463 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14608 7554 7463 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14607 3625 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14606 3625 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14605 8144 5648 3625 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14604 8144 3857 3625 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14603 3628 7026 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14602 3628 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14601 8144 6797 3628 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14600 8144 6544 3628 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14599 3865 4474 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14598 8144 4311 3865 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14597 3258 4292 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14596 8144 4468 3258 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14595 2680 2679 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14594 8144 5453 2680 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14593 2887 2680 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14592 2839 3759 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14591 8144 4166 2839 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14590 2836 2839 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14589 3136 4947 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14588 8144 3134 3136 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14587 3135 3136 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14586 2647 2868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14585 8144 3229 2647 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14584 2853 2647 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14583 6157 6906 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14582 8144 6905 6157 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14581 8144 713 710 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14580 713 939 602 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14579 603 714 713 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14578 8144 939 714 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14577 602 4160 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14576 8144 709 603 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14575 710 713 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14574 8144 548 549 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14573 548 939 461 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14572 460 462 548 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14571 8144 939 462 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14570 461 4176 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14569 8144 535 460 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14568 549 548 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14567 8144 294 292 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14566 294 939 228 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14565 227 296 294 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14564 8144 939 296 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14563 228 3999 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14562 8144 514 227 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14561 292 294 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14560 8144 322 320 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14559 322 939 232 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14558 231 324 322 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14557 8144 939 324 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14556 232 2402 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14555 8144 532 231 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14554 320 322 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14553 8144 2403 2402 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14552 2403 5148 2300 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14551 2299 2406 2403 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14550 8144 5148 2406 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14549 2300 8122 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14548 8144 6076 2299 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14547 2402 2403 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14546 1145 1996 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14545 1145 4540 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14544 8144 5148 1145 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14543 8144 1372 1145 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14542 5054 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14541 5139 5907 5054 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14540 8144 6549 5139 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14539 2941 2462 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14538 2941 2240 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14537 8144 2935 2941 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14536 1420 1761 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14535 1741 1760 1420 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14534 8144 3148 1741 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14533 7002 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14532 7002 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14531 8144 7356 7002 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14530 8144 6292 7002 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14529 8144 4173 3988 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14528 3988 4172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14527 8144 7349 3988 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14526 3987 3988 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14525 8144 5428 5425 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14524 5425 5424 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14523 8144 5619 5425 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14522 5911 5425 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14521 8144 4529 4528 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14520 4528 4548 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14519 8144 4527 4528 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14518 6294 4528 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14517 8144 672 671 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14516 672 903 592 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14515 591 675 672 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14514 8144 903 675 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14513 592 3537 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14512 8144 677 591 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14511 671 672 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14510 8144 3540 3537 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14509 3540 4178 3539 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14508 3538 3541 3540 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14507 8144 4178 3541 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14506 3539 4662 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14505 8144 7549 3538 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14504 3537 3540 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14503 8144 6992 6985 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14502 8144 7957 6986 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14501 6985 6986 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14500 8144 5654 4218 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14499 4218 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14498 4218 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14497 8144 5938 4218 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14496 4503 4218 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14495 7879 7876 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14494 7878 7877 7879 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14493 8144 7889 7878 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14492 3968 5938 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14491 3968 6520 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14490 8144 5453 3968 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14489 8144 5606 3968 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14488 4200 5150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14487 8144 4439 4200 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14486 4198 4200 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14485 3144 3146 3067 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14484 8144 4510 3067 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14483 3067 4007 3144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14482 3145 3144 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14481 8144 5898 5587 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14480 8144 8064 5404 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14479 5587 5404 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14478 6958 7296 6957 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14477 6957 7885 7128 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14476 7128 7877 6958 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14475 6958 7884 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14474 8144 7869 6958 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14473 7126 7128 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14472 5378 5383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14471 8144 6793 5378 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14470 5377 5378 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14469 3163 3170 3164 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14468 3164 3171 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14467 8144 4742 3163 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14466 3250 3163 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14465 3633 4071 3632 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14464 3630 3635 3633 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14463 3631 3629 3630 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14462 8144 3636 3631 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14461 3651 3632 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14460 1089 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14459 8144 1088 1089 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14458 1760 1089 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14457 1050 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14456 8144 1048 1050 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14455 1476 1050 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14454 5540 5669 5668 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14453 8144 7352 5669 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14452 5541 6359 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14451 5668 7352 5541 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14450 8144 6358 5540 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14449 8144 7888 7123 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14448 7123 7619 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14447 7123 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14446 8144 8184 7123 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14445 7121 7123 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14444 2225 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14443 2226 7343 2225 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14442 2224 4540 2226 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14441 8144 2698 2224 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14440 2234 2226 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14439 8144 6597 6601 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14438 6598 6594 6453 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14437 6453 6597 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14436 6453 6601 6598 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14435 8144 6596 6453 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14434 6596 6594 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14433 2881 4517 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14432 8144 4518 2881 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14431 4203 2881 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14430 2180 2178 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14429 2181 2179 2180 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14428 8144 4429 2181 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14427 554 7548 555 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14426 555 1798 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14425 8144 6363 554 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14424 557 554 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14423 2762 7779 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14422 2886 7778 2762 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14421 8144 8122 2886 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14420 7431 7559 7430 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14419 7430 7548 7539 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14418 7539 7550 7431 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14417 7431 8051 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14416 8144 8061 7431 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14415 7536 7539 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14414 8144 1565 1567 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14413 1567 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14412 8144 4306 1567 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14411 4178 1567 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14410 1727 2346 1728 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14409 1728 2610 1727 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14408 8144 2616 1728 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14407 4106 4939 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14406 4189 5406 4106 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14405 8144 6553 4189 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14404 5569 5633 5529 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14403 5529 5567 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14402 8144 6763 5569 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14401 5566 5569 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14400 8144 5648 2042 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14399 2042 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14398 2042 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14397 8144 5447 2042 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14396 2043 2042 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14395 8139 7612 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14394 7777 6988 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14393 8144 6396 5033 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14392 5033 5875 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14391 5033 6172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14390 8144 6921 5033 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14389 5032 5033 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14388 8144 6914 5734 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14387 5734 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14386 8144 7130 5734 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14385 5732 5734 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14384 221 1115 222 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14383 222 1114 271 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14382 271 273 222 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14381 221 266 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14380 8144 1110 221 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14379 222 268 221 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14378 1744 271 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14377 8144 2430 2209 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14376 2209 2424 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14375 2209 2421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14374 8144 4203 2209 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14373 2407 2209 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14372 4147 4416 4101 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14371 4101 4152 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14370 8144 4156 4147 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14369 4492 4147 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14368 128 129 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14367 124 130 123 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14366 8144 529 124 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14365 130 131 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14364 8144 1772 131 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14363 8144 306 129 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14362 126 130 128 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14361 127 131 126 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14360 8144 125 127 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14359 125 126 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14358 123 131 125 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14357 8144 123 529 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14356 529 123 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14355 4456 4561 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14354 4454 4562 4557 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14353 8144 4558 4454 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14352 4562 4563 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14351 8144 5864 4563 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14350 8144 4765 4561 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14349 4560 4562 4456 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14348 4455 4563 4560 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14347 8144 4559 4455 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14346 4559 4560 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14345 4557 4563 4559 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14344 8144 4557 4558 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14343 4558 4557 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14342 7535 7778 7429 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14341 7429 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14340 8144 7549 7535 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14339 7768 7535 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14338 1424 4025 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14337 1525 1778 1424 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14336 8144 4198 1525 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14335 2863 2875 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14334 8144 2873 2863 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14333 611 737 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14332 609 736 730 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14331 8144 1111 609 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14330 736 738 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14329 8144 1772 738 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14328 8144 920 737 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14327 732 736 611 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14326 610 738 732 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14325 8144 733 610 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14324 733 732 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14323 730 738 733 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14322 8144 730 1111 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14321 1111 730 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14320 7362 7778 7262 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14319 7262 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14318 8144 8139 7362 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14317 7357 7362 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14316 1530 5136 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14315 8144 1497 1530 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14314 7559 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14313 8144 7026 7559 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14312 4026 4024 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14311 7406 4025 4026 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14310 8144 4207 7406 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14309 6555 6835 6440 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14308 6440 8058 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14307 8144 6554 6555 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14306 6553 6555 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14305 2652 2868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14304 8144 3229 2652 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14303 7809 7811 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14302 7805 7812 7806 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14301 8144 8059 7805 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14300 7812 7813 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14299 8144 8063 7813 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14298 8144 8122 7811 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14297 7810 7812 7809 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14296 7808 7813 7810 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14295 8144 7807 7808 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14294 7807 7810 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14293 7806 7813 7807 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14292 8144 7806 8059 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14291 8059 7806 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14290 68 70 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14289 64 71 65 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14288 8144 6484 64 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14287 71 72 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14286 8144 1951 72 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14285 8144 3511 70 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14284 69 71 68 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14283 66 72 69 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14282 8144 67 66 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14281 67 69 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14280 65 72 67 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14279 8144 65 6484 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14278 6484 65 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14277 8144 3588 3596 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14276 3588 8064 3590 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14275 3589 3591 3588 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14274 8144 8064 3591 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14273 3590 3787 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14272 8144 4712 3589 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14271 3596 3588 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14270 6959 7158 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14269 7135 7877 6959 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14268 8144 7885 7135 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14267 6420 8187 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14266 6421 7893 6420 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14265 8144 7869 6421 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14264 3700 4798 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14263 3858 3856 3700 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14262 8144 3857 3858 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14261 531 1115 533 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14260 533 1114 534 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14259 534 532 533 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14258 531 529 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14257 8144 1110 531 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14256 533 530 531 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14255 2179 534 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14254 7327 8040 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14253 7327 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14252 8144 7352 7327 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14251 2206 2968 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14250 2206 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14249 8144 4572 2206 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14248 7286 7383 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14247 7284 7385 7378 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14246 8144 7379 7284 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14245 7385 7382 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14244 8144 8166 7382 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14243 8144 7384 7383 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14242 7381 7385 7286 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14241 7285 7382 7381 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14240 8144 7380 7285 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14239 7380 7381 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14238 7378 7382 7380 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14237 8144 7378 7379 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14236 7379 7378 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14235 6757 6759 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14234 6753 6760 6754 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14233 8144 7513 6753 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14232 6760 6761 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14231 8144 8063 6761 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_14230 8144 7485 6759 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14229 6758 6760 6757 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14228 6756 6761 6758 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14227 8144 6755 6756 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14226 6755 6758 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14225 6754 6761 6755 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_14224 8144 6754 7513 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14223 7513 6754 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14222 8144 2194 2398 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14221 2194 8094 2195 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14220 2193 2196 2194 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14219 8144 8094 2196 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14218 2195 2390 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14217 8144 6080 2193 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14216 2398 2194 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14215 8144 3092 3282 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14214 3092 8094 3064 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14213 3062 3065 3092 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14212 8144 8094 3065 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14211 3064 3063 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14210 8144 5563 3062 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14209 3282 3092 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14208 8144 3298 3519 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14207 3298 8094 3202 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14206 3201 3301 3298 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14205 8144 8094 3301 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14204 3202 3300 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14203 8144 5387 3201 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14202 3519 3298 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14201 8144 1309 1307 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14200 1309 8094 1308 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14199 1310 1311 1309 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14198 8144 8094 1311 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14197 1308 1474 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14196 8144 5394 1310 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14195 1307 1309 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14194 8144 1521 1519 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14193 1521 8094 1423 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14192 1422 1523 1521 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14191 8144 8094 1523 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14190 1423 1525 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14189 8144 5419 1422 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14188 1519 1521 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14187 8144 1492 1488 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14186 1492 8094 1418 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14185 1417 1493 1492 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14184 8144 8094 1493 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14183 1418 1490 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14182 8144 5571 1417 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14181 1488 1492 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14180 5114 5606 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14179 5114 5108 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14178 8144 5938 5114 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14177 3300 2805 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14176 8144 1052 3300 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14175 764 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14174 8144 5483 764 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14173 1945 3348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14172 8144 3315 1945 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14171 2616 1945 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14170 1920 2796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14169 8144 3542 1920 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14168 2135 1920 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14167 3777 3780 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14166 8144 4543 3777 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14165 3774 3777 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14164 3543 3586 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14163 3543 3989 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14162 8144 3990 3543 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14161 8144 3581 3543 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14160 2657 2877 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14159 2661 2866 2657 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14158 8144 7314 2661 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14157 8144 1979 1974 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14156 1979 8094 1853 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14155 1852 1980 1979 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14154 8144 8094 1980 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14153 1853 1978 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14152 8144 5435 1852 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14151 1974 1979 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14150 8144 1529 1526 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14149 1529 8094 1426 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14148 1425 1531 1529 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14147 8144 8094 1531 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14146 1426 1530 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14145 8144 5443 1425 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14144 1526 1529 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14143 8144 1970 2189 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14142 1970 8094 1851 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14141 1850 1972 1970 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14140 8144 8094 1972 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14139 1851 2182 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14138 8144 5143 1850 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_14137 2189 1970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14136 4725 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14135 4725 7354 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14134 8144 4572 4725 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14133 8144 6143 4725 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14132 3199 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14131 4129 5907 3199 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14130 8144 6292 4129 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14129 1421 1760 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14128 1497 1761 1421 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14127 8144 8045 1497 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14126 2946 4470 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14125 8144 3033 2946 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14124 1696 2698 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14123 1802 1887 1696 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14122 1695 1986 1802 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14121 8144 2926 1695 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14120 3253 1802 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14119 3608 5483 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14118 3608 4051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14117 8144 4572 3608 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14116 1148 774 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14115 1148 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14114 8144 4572 1148 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14113 1553 2687 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14112 1553 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14111 8144 6543 1553 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14110 8144 7327 7326 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14109 7326 7328 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14108 8144 7329 7326 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14107 7325 7326 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14106 8144 3759 3113 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14105 3113 4166 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14104 8144 3744 3113 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14103 3111 3113 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14102 8144 3763 3125 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14101 3125 4424 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14100 8144 3744 3125 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14099 3123 3125 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14098 1792 1362 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14097 1792 1361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14096 8144 1550 1792 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14095 8144 1553 1792 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14094 2439 2693 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14093 2439 2441 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14092 8144 2437 2439 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14091 8144 2913 2439 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14090 6822 6821 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14089 6820 7058 6822 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14088 8144 7053 6820 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14087 1432 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14086 1580 1891 1432 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14085 1431 1996 1580 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14084 8144 2698 1431 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14083 2233 1580 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14082 2723 4167 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14081 2723 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14080 8144 6797 2723 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14079 8144 4306 2723 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14078 5265 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14077 5265 6396 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14076 8144 6172 5265 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14075 8144 6921 5265 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14074 8144 2254 1871 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14073 1871 2252 2031 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14072 2032 2031 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14071 4320 5041 4116 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14070 4116 4583 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14069 8144 4317 4320 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14068 4318 4320 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14067 6431 6502 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14066 6513 6503 6431 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14065 8144 6504 6513 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14064 6916 7305 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14063 6915 7301 6916 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14062 8144 6914 6915 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14061 2776 2926 2920 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14060 2775 3170 2776 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14059 8144 3171 2775 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14058 2919 2920 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14057 5534 6090 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14056 5900 6089 5534 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14055 8144 6576 5900 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14054 4166 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14053 4166 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14052 8144 4167 4166 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14051 8144 6506 4166 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14050 8144 7403 7402 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14049 7402 7884 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14048 8144 7883 7402 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14047 8179 7402 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14046 3672 3716 3715 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14045 3673 7787 3672 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14044 3671 8048 3673 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14043 8144 8045 3671 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_14042 3714 3715 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14041 4138 4898 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14040 8144 4405 4138 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14039 4137 4138 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14038 1551 1559 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14037 8144 2924 1551 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14036 1550 1551 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14035 2455 2469 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14034 8144 4572 2455 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14033 2707 2455 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14032 2218 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14031 8144 4574 2218 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14030 2896 2218 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14029 1045 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14028 8144 1043 1045 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14027 1743 1045 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14026 6789 6835 6790 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14025 6790 7280 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14024 8144 7025 6789 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14023 6788 6789 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14022 4019 7791 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14021 4018 7788 4019 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14020 8144 6080 4018 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14019 5382 5633 5381 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14018 5381 5380 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14017 8144 5817 5382 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14016 5379 5382 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14015 5423 5633 5422 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14014 5422 5421 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14013 8144 7536 5423 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14012 5420 5423 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_14011 5975 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14010 8144 8184 5975 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14009 5879 5975 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14008 8144 359 164 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14007 164 1150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14006 8144 3384 164 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_14005 163 164 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14004 8144 3744 3680 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14003 3680 3991 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14002 4143 3740 3680 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14001 3679 3737 4143 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_14000 3680 4141 3679 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13999 5928 6019 5848 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13998 5848 5929 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13997 8144 5927 5928 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13996 6102 5928 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13995 8144 2454 2250 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13994 2250 2249 2251 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13993 8144 5041 5043 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13992 5043 5273 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13991 5043 5269 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13990 8144 5042 5043 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13989 5040 5043 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13988 7248 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13987 7323 7798 7248 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13986 8144 7585 7323 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13985 2266 2269 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13984 2263 2270 2264 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13983 8144 2262 2263 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13982 2270 2271 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13981 8144 3834 2271 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13980 8144 3193 2269 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13979 2267 2270 2266 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13978 2268 2271 2267 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13977 8144 2265 2268 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13976 2265 2267 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13975 2264 2271 2265 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13974 8144 2264 2262 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13973 2262 2264 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13972 5068 5209 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13971 5066 5210 5204 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13970 8144 5202 5066 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13969 5210 5211 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13968 8144 5864 5211 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13967 8144 5487 5209 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13966 5207 5210 5068 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13965 5067 5211 5207 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13964 8144 5205 5067 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13963 5205 5207 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13962 5204 5211 5205 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13961 8144 5204 5202 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13960 5202 5204 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13959 4313 4583 4114 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13958 4114 5265 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13957 8144 4312 4313 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13956 4311 4313 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13955 8144 5940 2030 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13954 2030 2262 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13953 2030 2964 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13952 8144 2968 2030 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13951 2469 2030 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13950 8144 1898 1820 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13949 1820 1897 2027 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13948 8144 4573 968 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13947 968 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13946 968 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13945 8144 4302 968 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13944 1618 968 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13943 8144 6797 3640 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13942 3640 3639 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13941 3640 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13940 8144 6293 3640 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13939 3856 3640 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13938 3132 3141 3131 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13937 3131 3552 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13936 8144 3553 3132 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13935 3130 3132 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13934 3277 3964 3198 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13933 3198 3276 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13932 8144 4503 3277 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13931 3275 3277 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13930 151 152 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13929 147 153 146 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13928 8144 532 147 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13927 153 154 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13926 8144 3834 154 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13925 8144 320 152 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13924 149 153 151 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13923 150 154 149 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13922 8144 148 150 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13921 148 149 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13920 146 154 148 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13919 8144 146 532 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13918 532 146 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13917 942 565 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13916 942 557 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13915 8144 763 942 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13914 1535 1539 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13913 1535 1782 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13912 8144 4172 1535 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13911 1541 1539 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13910 1541 1538 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13909 8144 4172 1541 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13908 3193 3191 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13907 8144 3192 3193 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13906 4020 4021 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13905 4208 7788 4020 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13904 8144 6541 4208 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13903 3958 5099 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13902 8144 1466 3958 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13901 3353 3150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13900 8144 6363 3353 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13899 4950 5406 4949 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13898 4949 7059 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13897 8144 6834 4950 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13896 4947 4950 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13895 4972 4974 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13894 4968 4975 4969 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13893 8144 5180 4968 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13892 4975 4976 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13891 8144 5864 4976 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13890 8144 5181 4974 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13889 4973 4975 4972 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13888 4971 4976 4973 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13887 8144 4970 4971 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13886 4970 4973 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13885 4969 4976 4970 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13884 8144 4969 5180 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13883 5180 4969 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13882 1401 1484 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13881 1399 1486 1479 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13880 8144 5571 1399 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13879 1486 1487 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13878 8144 1951 1487 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13877 8144 1488 1484 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13876 1483 1486 1401 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13875 1400 1487 1483 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13874 8144 1481 1400 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13873 1481 1483 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13872 1479 1487 1481 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13871 8144 1479 5571 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13870 5571 1479 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13869 4499 4668 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13868 4493 4615 4665 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13867 8144 5108 4493 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13866 4615 4669 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13865 8144 8063 4669 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13864 8144 4666 4668 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13863 4614 4615 4499 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13862 4496 4669 4614 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13861 8144 4612 4496 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13860 4612 4614 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13859 4665 4669 4612 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13858 8144 4665 5108 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13857 5108 4665 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13856 7751 7766 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13855 7749 7747 7751 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13854 8144 7748 7749 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13853 5415 5413 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13852 5414 5432 5415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13851 8144 5436 5414 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13850 8175 7890 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13849 8144 7887 8175 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13848 7875 7878 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13847 8144 7874 7875 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13846 7399 6915 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13845 8144 6912 7399 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13844 6627 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13843 8144 6618 6627 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13842 3853 3867 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13841 8144 4292 3853 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13840 2169 4171 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13839 2630 2167 2169 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13838 8144 2375 2630 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13837 3090 3284 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13836 3082 3283 3279 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13835 8144 5563 3082 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13834 3283 3285 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13833 8144 3708 3285 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13832 8144 3282 3284 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13831 3227 3283 3090 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13830 3087 3285 3227 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13829 8144 3226 3087 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13828 3226 3227 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13827 3279 3285 3226 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13826 8144 3279 5563 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13825 5563 3279 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13824 7031 7053 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13823 8144 7343 7031 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13822 7339 7031 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13821 7034 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13820 7034 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13819 8144 7356 7034 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13818 8144 6349 7034 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13817 6897 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13816 8144 6883 6897 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13815 5501 6412 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13814 5501 5500 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13813 8144 6415 5501 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13812 1806 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13811 1806 7026 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13810 8144 5654 1806 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13809 7149 7408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13808 8144 8184 7149 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13807 8144 6343 6590 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13806 6343 6838 6345 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13805 6342 6346 6343 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13804 8144 6838 6346 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13803 6345 6344 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13802 8144 6341 6342 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13801 6590 6343 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13800 8144 6592 6597 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13799 6592 6864 6452 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13798 6451 6593 6592 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13797 8144 6864 6593 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13796 6452 6590 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13795 8144 6588 6451 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13794 6597 6592 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13793 3661 3660 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13792 8144 4074 3661 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13791 8144 6090 4948 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13790 4946 4948 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13789 8144 7343 4946 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13788 4945 4946 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13787 8144 4946 4945 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13786 4943 5147 4944 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13785 8144 7955 4944 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13784 4944 5148 4943 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13783 4942 4943 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13782 2345 3097 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13781 8144 3553 2345 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13780 2344 2345 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13779 3117 3316 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13778 8144 3229 3117 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13777 3559 3117 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13776 3763 7863 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13775 3763 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13774 8144 4172 3763 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13773 8144 94 91 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13772 94 903 92 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13771 93 95 94 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13770 8144 903 95 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13769 92 3532 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13768 8144 268 93 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13767 91 94 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13766 7012 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13765 7012 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13764 8144 7026 7012 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13763 8144 8000 7012 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13762 1001 1476 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13761 1047 1477 1001 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13760 8144 8045 1047 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13759 1891 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13758 1891 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13757 8144 4306 1891 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13756 5871 7893 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13755 5968 7408 5871 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13754 8144 8184 5968 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13753 5269 6172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13752 5269 5875 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13751 8144 6396 5269 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13750 8144 6672 5269 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13749 8144 6568 6588 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13748 6568 6838 6445 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13747 6444 6571 6568 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13746 8144 6838 6571 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13745 6445 6823 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13744 8144 6567 6444 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13743 6588 6568 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13742 3867 4061 3697 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13741 3697 3841 3867 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13740 8144 4280 3697 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13739 1812 1996 1811 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13738 1811 2926 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13737 8144 1813 1812 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13736 2239 1812 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13735 2430 2968 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13734 2430 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13733 8144 4293 2430 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13732 1999 5940 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13731 1999 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13730 8144 5483 1999 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13729 7742 7738 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13728 7742 7734 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13727 8144 7729 7742 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13726 8144 7730 7742 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13725 8144 3535 3532 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13724 3535 4178 3534 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13723 3533 3536 3535 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13722 8144 4178 3536 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13721 3534 4403 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13720 8144 7528 3533 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13719 3532 3535 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13718 6794 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13717 6794 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13716 8144 7026 6794 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13715 8144 8021 6794 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13714 3618 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13713 3618 3639 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13712 8144 7356 3618 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13711 8144 6293 3618 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13710 7006 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13709 7006 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13708 8144 6797 7006 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13707 8144 6520 7006 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13706 8144 3608 3366 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13705 3366 5168 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13704 8144 3373 3366 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13703 3610 3366 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13702 1722 2813 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_13701 1724 1719 1720 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13700 1720 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13699 8144 1721 1725 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13698 1725 1727 1723 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13697 1723 1722 1724 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13696 1724 2813 1726 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13695 1726 2610 1725 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13694 8144 3556 1721 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_13693 2589 1724 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13692 8144 4143 3985 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13691 4149 3986 3984 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13690 3984 4143 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13689 3984 3985 4149 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13688 8144 3983 3984 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13687 3983 3986 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13686 8144 264 261 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13685 264 903 220 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13684 219 265 264 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13683 8144 903 265 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13682 220 3978 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13681 8144 498 219 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13680 261 264 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13679 4593 4715 6850 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13678 8144 7314 4715 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13677 4594 4714 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13676 6850 7314 4594 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13675 8144 4712 4593 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13674 5122 5121 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13673 8144 5606 5122 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13672 5120 5122 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13671 5920 6127 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13670 8144 6576 5920 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13669 5846 5920 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13668 5899 6288 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13667 8144 5900 5899 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13666 5828 5899 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13665 7762 7760 7763 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13664 7763 7761 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13663 8144 7979 7762 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13662 7759 7762 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13661 5100 5406 5050 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13660 5050 6524 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13659 8144 5124 5100 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13658 5099 5100 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13657 8144 1924 246 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13656 1287 1711 216 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13655 216 1924 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13654 216 246 1287 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13653 8144 244 216 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13652 244 1711 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13651 8144 6541 3971 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13650 8144 8064 3973 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13649 3971 3973 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13648 646 2315 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13647 8144 3078 646 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13646 2806 646 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13645 2717 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13644 8144 4572 2717 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13643 2937 2717 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13642 1814 2027 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13641 8144 2235 1814 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13640 1817 1814 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13639 8144 6484 3765 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13638 8144 8064 3767 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13637 3765 3767 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13636 6044 6050 5977 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13635 8144 6274 5977 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13634 5977 6262 6044 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13633 6043 6044 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13632 6430 6500 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13631 6781 6783 6430 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13630 8144 7314 6781 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13629 8144 5453 4486 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13628 4486 5938 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13627 8144 5606 4486 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13626 4402 4486 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13625 6633 7881 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13624 8144 7891 6633 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13623 6632 6633 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13622 8144 8187 5972 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13621 5972 7893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13620 8144 7883 5972 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13619 5875 5972 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13618 5510 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13617 8144 7130 5510 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13616 6912 5510 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13615 8144 4302 953 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13614 953 5483 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13613 8144 5940 953 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13612 1133 953 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13611 1429 1546 5620 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13610 1428 1547 1429 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13609 8144 1545 1428 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13608 6333 6332 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13607 6331 6340 6333 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13606 6330 6334 6331 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13605 8144 7788 6330 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13604 6329 6331 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13603 5213 5695 5069 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13602 5069 5869 5213 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13601 8144 5212 5069 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13600 7863 7591 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13599 8122 8058 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13598 8144 6609 3824 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13597 3824 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13596 8144 5654 3824 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13595 7788 3824 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13594 8144 2951 2783 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13593 2783 2950 3877 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13592 2711 2706 2708 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13591 2708 2707 2709 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13590 2709 4295 2711 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13589 2711 5492 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13588 8144 4790 2711 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13587 2705 2709 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13586 8144 1543 1152 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13585 1152 1154 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13584 1152 1559 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13583 8144 1806 1152 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13582 1150 1152 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13581 870 873 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13580 867 874 868 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13579 8144 1048 867 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13578 874 875 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13577 8144 1951 875 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13576 8144 890 873 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13575 871 874 870 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13574 872 875 871 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13573 8144 869 872 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13572 869 871 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13571 868 875 869 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13570 8144 868 1048 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13569 1048 868 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13568 7366 7788 7266 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13567 7266 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13566 8144 8097 7366 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13565 7368 7366 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13564 7112 7379 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13563 234 354 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13562 335 334 234 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13561 233 342 335 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13560 8144 343 233 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13559 1110 335 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13558 4158 4157 4103 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13557 4103 4498 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13556 8144 4155 4158 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13555 4156 4158 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13554 3155 3386 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13553 3153 3387 3382 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13552 8144 3384 3153 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13551 3387 3388 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13550 8144 3834 3388 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13549 8144 4757 3386 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13548 3242 3387 3155 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13547 3154 3388 3242 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13546 8144 3241 3154 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13545 3241 3242 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13544 3382 3388 3241 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13543 8144 3382 3384 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13542 3384 3382 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13541 5424 6480 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13540 8144 5603 5424 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13539 3141 3146 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13538 8144 4007 3141 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13537 109 111 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13536 105 112 106 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13535 8144 703 105 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13534 112 113 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13533 8144 1951 113 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13532 8144 697 111 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13531 110 112 109 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13530 108 113 110 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13529 8144 107 108 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13528 107 110 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13527 106 113 107 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13526 8144 106 703 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13525 703 106 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13524 978 1036 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13523 976 1035 1030 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13522 8144 6267 976 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13521 1035 1037 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13520 8144 3708 1037 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13519 8144 6085 1036 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13518 1033 1035 978 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13517 977 1037 1033 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13516 8144 1031 977 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13515 1031 1033 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13514 1030 1037 1031 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13513 8144 1030 6267 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13512 6267 1030 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13511 8144 5661 5658 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13510 5661 6358 5521 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13509 5520 5662 5661 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13508 8144 6358 5662 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13507 5521 6076 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13506 8144 6142 5520 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13505 5658 5661 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13504 2182 4693 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13503 8144 2181 2182 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13502 2702 3158 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13501 8144 3857 2702 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13500 3129 3768 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13499 8144 3128 3129 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13498 7295 7393 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13497 7293 7389 7388 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13496 8144 7604 7293 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13495 7389 7390 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13494 8144 8166 7390 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13493 8144 7603 7393 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13492 7392 7389 7295 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13491 7294 7390 7392 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13490 8144 7391 7294 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13489 7391 7392 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13488 7388 7390 7391 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13487 8144 7388 7604 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13486 7604 7388 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13485 1138 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13484 8144 1372 1138 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13483 1359 1138 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13482 8144 4273 4271 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13481 4273 7871 4097 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13480 4098 4275 4273 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13479 8144 7871 4275 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13478 4097 4788 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13477 8144 4270 4098 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13476 4271 4273 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13475 5118 6549 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13474 5118 5121 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13473 8144 5606 5118 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13472 4795 5740 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13471 4795 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13470 8144 7887 4795 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13469 6004 6189 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13468 6186 7299 6004 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13467 6003 6667 6186 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13466 8144 6188 6003 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13465 6185 6186 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13464 4202 6089 4017 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13463 4017 4029 4202 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13462 8144 6090 4017 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13461 3780 3373 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13460 3780 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13459 8144 5168 3780 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13458 5171 5169 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13457 8144 5168 5171 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13456 6835 5171 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13455 6925 6970 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13454 6923 6969 6964 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13453 8144 7247 6923 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13452 6969 6971 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13451 8144 8063 6971 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13450 8144 7241 6970 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13449 6967 6969 6925 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13448 6924 6971 6967 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13447 8144 6965 6924 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13446 6965 6967 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13445 6964 6971 6965 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13444 8144 6964 7247 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13443 7247 6964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13442 7046 7062 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13441 8144 7343 7046 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13440 7543 7046 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13439 5079 5078 5045 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13438 5045 6477 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13437 8144 7957 5079 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13436 5077 5079 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13435 5044 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13434 8144 7130 5044 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13433 3623 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13432 3623 3826 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13431 8144 7356 3623 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13430 8144 5942 3623 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13429 4048 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13428 4048 4047 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13427 8144 6311 4048 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13426 8144 6293 4048 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13425 8144 1799 381 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13424 379 381 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13423 8144 2492 379 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13422 378 379 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13421 8144 379 378 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13420 2306 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13419 2452 4517 2306 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13418 2305 7343 2452 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13417 8144 2698 2305 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13416 2448 2452 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13415 5992 6090 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13414 6302 6089 5992 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13413 8144 6823 6302 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13412 7509 7508 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13411 8144 7512 7509 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13410 7753 7509 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13409 3990 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13408 3990 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13407 8144 4574 3990 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13406 8144 6775 3990 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13405 8144 2164 2166 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13404 2164 3114 2163 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13403 2161 2162 2164 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13402 8144 3114 2162 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13401 2163 3348 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13400 8144 3315 2161 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13399 2166 2164 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13398 5895 5896 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13397 8144 7343 5895 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13396 5825 5895 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13395 2906 3379 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13394 2906 4517 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13393 8144 3378 2906 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13392 8144 5169 2906 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13391 8144 4576 4570 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13390 4576 7871 4467 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13389 4465 4466 4576 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13388 8144 7871 4466 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13387 4467 6648 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13386 8144 4734 4465 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13385 4570 4576 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13384 5488 6629 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13383 5487 5494 5488 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13382 8144 5486 5487 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13381 8144 2492 374 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13380 372 374 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13379 8144 1799 372 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13378 375 372 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13377 8144 372 375 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13376 3072 3371 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13375 3152 3370 3072 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13374 3071 4302 3152 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13373 8144 5624 3071 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13372 7797 3152 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13371 955 5147 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13370 955 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13369 8144 1154 955 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13368 8144 1543 955 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13367 8144 7088 7398 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13366 7088 7867 6938 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13365 6937 7090 7088 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13364 8144 7867 7090 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13363 6938 7528 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13362 8144 7572 6937 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13361 7398 7088 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13360 4204 4203 4107 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13359 4107 4705 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13358 8144 4202 4204 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13357 4206 4204 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13356 8144 2421 2417 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13355 2417 2430 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13354 2417 4203 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13353 8144 2924 2417 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13352 5406 2417 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13351 8144 4901 4903 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13350 4903 4902 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13349 8144 5606 4903 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13348 4900 4903 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13347 4583 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13346 4583 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13345 8144 5483 4583 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13344 8144 4075 4583 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13343 4301 4473 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13342 8144 4298 4301 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13341 4299 4301 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13340 4516 5399 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13339 8144 4956 4516 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13338 4437 4516 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13337 593 1115 594 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13336 594 1114 681 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13335 681 1063 594 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13334 593 676 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13333 8144 1110 593 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13332 594 677 593 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13331 1477 681 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13330 2158 2822 2157 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13329 2157 2156 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13328 8144 3315 2158 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13327 2155 2158 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13326 1847 1964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13325 2177 1965 1847 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13324 8144 1962 2177 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13323 8144 3570 3323 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13322 3577 3567 3208 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13321 3208 3570 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13320 3208 3323 3577 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13319 8144 3324 3208 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13318 3324 3567 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13317 8144 6489 6279 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13316 8144 7500 6277 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13315 6279 6277 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13314 5385 5384 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13313 8144 5606 5385 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13312 5390 5385 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13311 8144 7026 1378 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13310 1378 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13309 1378 4572 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13308 8144 5447 1378 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13307 1377 1378 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13306 8144 5648 3389 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13305 3389 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13304 3389 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13303 8144 3857 3389 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13302 3390 3389 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13301 8144 4068 3369 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13300 3369 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13299 8144 4293 3369 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13298 4021 3369 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13297 2751 2975 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13296 2749 2976 2970 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13295 8144 2968 2749 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13294 2976 2977 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13293 8144 3834 2977 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13292 8144 3197 2975 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13291 2972 2976 2751 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13290 2750 2977 2972 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13289 8144 2971 2750 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13288 2971 2972 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13287 2970 2977 2971 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13286 8144 2970 2968 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13285 2968 2970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13284 8144 8064 467 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13283 466 467 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13282 8144 3077 466 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13281 1909 466 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13280 8144 466 1909 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13279 6815 7778 6817 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13278 6817 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13277 8144 7349 6815 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13276 6816 6815 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13275 8144 4468 2952 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13274 2952 2955 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13273 2952 2958 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13272 8144 2957 2952 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13271 3186 2952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13270 2697 2696 2917 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13269 2694 2904 2697 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13268 8144 2695 2694 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13267 2772 2919 3167 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13266 2771 2917 2772 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13265 8144 3251 2771 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13264 8144 3644 3189 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13263 3188 3189 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13262 8144 3187 3188 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13261 3191 3188 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13260 8144 3188 3191 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13259 8144 2723 2475 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13258 2475 2722 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13257 2475 2481 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13256 8144 2473 2475 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13255 2471 2475 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13254 6943 7103 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13253 6941 7102 7097 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13252 8144 7095 6941 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13251 7102 7105 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13250 8144 8166 7105 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13249 8144 7108 7103 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13248 7101 7102 6943 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13247 6942 7105 7101 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13246 8144 7098 6942 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13245 7098 7101 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13244 7097 7105 7098 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13243 8144 7097 7095 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13242 7095 7097 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13241 4941 6294 4940 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13240 4940 4939 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13239 8144 5144 4941 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13238 5428 4941 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13237 8144 2439 1857 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13236 1858 2216 1890 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13235 1859 2005 1858 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13234 1857 1889 1859 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13233 2304 2682 2303 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13232 2441 7353 2304 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13231 2304 3371 2441 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13230 2303 4302 2304 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13229 2303 2896 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13228 8144 4306 2303 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13227 6836 6835 6837 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13226 6837 7591 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13225 8144 7062 6836 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13224 6834 6836 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13223 1410 1626 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13222 1408 1627 1621 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13221 8144 1799 1408 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13220 1627 1628 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13219 8144 3834 1628 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13218 8144 2961 1626 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13217 1623 1627 1410 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13216 1409 1628 1623 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13215 8144 1622 1409 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13214 1622 1623 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13213 1621 1628 1622 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13212 8144 1621 1799 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13211 1799 1621 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13210 1771 1770 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13209 1765 1773 1766 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13208 8144 5435 1765 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13207 1773 1774 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13206 8144 1772 1774 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13205 8144 1974 1770 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13204 1768 1773 1771 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13203 1769 1774 1768 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13202 8144 1767 1769 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13201 1767 1768 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13200 1766 1774 1767 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13199 8144 1766 5435 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13198 5435 1766 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13197 2275 2328 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13196 2273 2327 2322 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13195 8144 6292 2273 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13194 2327 2329 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13193 8144 3708 2329 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13192 8144 4641 2328 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13191 2325 2327 2275 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13190 2274 2329 2325 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13189 8144 2324 2274 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13188 2324 2325 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13187 2322 2329 2324 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13186 8144 2322 6292 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13185 6292 2322 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13184 946 1157 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13183 946 778 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13182 8144 1543 946 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13181 3373 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13180 3373 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13179 8144 5654 3373 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13178 4581 5038 4478 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13177 4478 4583 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13176 8144 4582 4581 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13175 4477 4581 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13174 4511 7777 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13173 4511 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13172 8144 4172 4511 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13171 923 1123 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13170 8144 1110 923 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13169 6955 7559 6954 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13168 6954 7548 7070 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13167 7070 7550 6955 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13166 6955 7263 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13165 8144 7264 6955 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13164 7068 7070 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13163 1157 5483 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13162 1157 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13161 8144 5654 1157 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13160 3244 3390 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13159 8144 6598 3244 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13158 8144 3583 3585 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13157 3584 3585 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13156 8144 3776 3584 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13155 3582 3584 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13154 8144 3584 3582 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13153 5400 6506 5398 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13152 5399 7247 5400 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13151 5400 6285 5399 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13150 5398 6286 5400 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13149 5398 6801 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13148 8144 6284 5398 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13147 3518 3520 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13146 3513 3521 3514 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13145 8144 5387 3513 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13144 3521 3522 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13143 8144 3708 3522 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_13142 8144 3519 3520 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13141 3517 3521 3518 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13140 3516 3522 3517 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13139 8144 3515 3516 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13138 3515 3517 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13137 3514 3522 3515 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13136 8144 3514 5387 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13135 5387 3514 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13134 7333 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13133 7333 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13132 8144 7356 7333 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13131 8144 6801 7333 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13130 5622 5620 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13129 8144 5618 5622 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13128 5619 5622 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13127 5718 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13126 5718 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13125 8144 6900 5718 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13124 2462 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13123 2462 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13122 8144 2469 2462 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13121 8144 2951 2309 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13120 2309 2950 2479 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13119 2477 2479 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13118 2202 1986 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13117 2202 2203 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13116 8144 5148 2202 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13115 7317 7747 7244 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13114 7244 7955 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13113 8144 7319 7317 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13112 7489 7317 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_13111 2147 2813 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_13110 2149 2144 2146 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13109 2146 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13108 8144 2145 2151 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13107 2151 2337 2148 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13106 2148 2147 2149 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13105 2149 2813 2150 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13104 2150 2340 2151 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13103 8144 3556 2145 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_13102 2143 2149 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13101 4990 4997 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_13100 4992 7612 4989 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13099 4989 6359 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13098 8144 4988 4994 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13097 4994 5202 4991 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13096 4991 4990 4992 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13095 4992 4997 4993 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13094 4993 7056 4994 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_13093 8144 6359 4988 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_13092 4987 4992 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13091 8144 3979 3978 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13090 3979 4178 3981 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13089 3980 3982 3979 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13088 8144 4178 3982 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13087 3981 5391 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13086 8144 7585 3980 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13085 3978 3979 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13084 7025 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13083 7025 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13082 8144 7026 7025 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13081 8144 8040 7025 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13080 4507 4712 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13079 8144 7314 4507 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13078 4286 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13077 4286 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13076 8144 7354 4286 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13075 8144 5654 4286 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13074 5031 5868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13073 5031 6636 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13072 8144 6921 5031 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13071 8144 7130 5031 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13070 4792 7887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13069 4792 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13068 8144 4790 4792 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13067 8144 7149 4792 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13066 8144 4143 4146 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13065 4497 4141 4100 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13064 4100 4143 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13063 4100 4146 4497 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13062 8144 4144 4100 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13061 4144 4141 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13060 2842 3759 2740 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13059 8144 4510 2740 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13058 2740 4166 2842 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13057 2840 2842 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13056 8144 550 751 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13055 550 903 464 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13054 463 465 550 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13053 8144 903 465 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13052 464 4012 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13051 8144 1116 463 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13050 751 550 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13049 8144 4014 4012 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13048 4014 5148 4013 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13047 4015 4016 4014 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13046 8144 5148 4016 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13045 4013 7349 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13044 8144 6541 4015 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13043 4012 4014 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13042 8144 901 899 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13041 901 903 904 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13040 902 905 901 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13039 8144 903 905 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13038 904 4160 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13037 8144 900 902 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13036 899 901 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13035 8144 4162 4160 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13034 4162 4178 4085 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13033 4084 4164 4162 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13032 8144 4178 4164 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13031 4085 4414 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13030 8144 7777 4084 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13029 4160 4162 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13028 4187 5837 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13027 8144 4428 4187 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13026 4184 4187 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13025 5411 5413 5412 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13024 5409 7787 5411 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13023 5410 8048 5409 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13022 8144 8045 5410 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13021 5408 5412 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13020 6946 6991 6988 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13019 8144 7957 6991 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_13018 6947 6992 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13017 6988 7957 6947 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13016 8144 6987 6946 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13015 1611 7026 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13014 1611 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13013 8144 4068 1611 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13012 8144 6796 1611 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_13011 3647 3851 3649 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13010 3648 3853 3647 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13009 3646 3645 3648 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13008 8144 3651 3646 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13007 3644 3649 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13006 2308 2466 2468 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13005 2307 2467 2308 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13004 8144 2705 2307 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_13003 2962 2468 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13002 7417 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13001 7512 7798 7417 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_13000 8144 7549 7512 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12999 8144 1924 866 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12998 865 2136 864 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12997 864 1924 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12996 864 866 865 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12995 8144 863 864 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12994 863 2136 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12993 8144 965 966 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12992 6802 966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12991 8144 966 6802 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12990 8144 966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12989 8144 966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12988 8144 965 784 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12987 6311 784 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12986 8144 784 6311 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12985 8144 784 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12984 8144 784 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12983 8144 574 572 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12982 965 572 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12981 8144 572 965 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12980 8144 572 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12979 8144 572 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12978 8144 7314 6275 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12977 6276 6275 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12976 8144 6273 6276 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12975 6274 6276 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12974 8144 6276 6274 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12973 780 2492 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12972 8144 1799 780 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12971 2718 780 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12970 4780 4782 4610 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12969 4610 5720 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12968 8144 7352 4780 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12967 4779 4780 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12966 3849 3847 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12965 8144 4792 3849 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12964 3850 3849 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12963 7396 7877 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12962 8144 7885 7396 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12961 7299 7396 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12960 3666 3868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12959 8144 3860 3666 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12958 3665 3666 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12957 5602 6062 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12956 8144 5838 5602 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12955 5600 5602 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12954 8144 7645 6922 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12953 6921 6922 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12952 8144 6922 6921 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12951 8144 6922 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12950 8144 6922 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12949 8144 7645 6673 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12948 6672 6673 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12947 8144 6673 6672 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12946 8144 6673 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12945 8144 6673 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12944 8144 7646 7647 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12943 7645 7647 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12942 8144 7647 7645 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12941 8144 7647 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12940 8144 7647 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12939 8144 7881 7153 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12938 7153 7403 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12937 7153 7884 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12936 8144 8184 7153 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12935 7405 7153 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12934 8144 7888 7141 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12933 7141 7643 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12932 7141 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12931 8144 7883 7141 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12930 7140 7141 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12929 8144 4018 2416 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12928 2416 2678 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12927 8144 2412 2416 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12926 2413 2416 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12925 2902 2901 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12924 8144 5908 2902 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12923 2912 2902 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12922 4732 4730 4599 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12921 4599 4955 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12920 8144 4731 4732 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12919 5680 4732 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12918 8144 760 556 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12917 556 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12916 8144 1891 556 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12915 559 556 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12914 5396 5406 5397 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12913 5397 6793 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12912 8144 6517 5396 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12911 5395 5396 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12910 8144 4575 2463 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12909 2463 2469 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12908 8144 4302 2463 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12907 2710 2463 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12906 7119 7604 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12905 8137 8147 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12904 7596 8125 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12903 5544 6629 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12902 5704 5710 5544 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12901 8144 5862 5704 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12900 7858 8119 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12899 5025 5015 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12898 4635 4558 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12897 3391 4270 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12896 4251 3384 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12895 5000 5485 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12894 8144 1893 1815 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12893 1815 2039 1818 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12892 2153 2156 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12891 2154 2822 2153 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12890 8144 3315 2154 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12889 2379 4003 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12888 8144 2177 2379 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12887 3329 3327 3209 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12886 3209 3552 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12885 8144 3553 3329 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12884 3569 3329 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12883 3682 3750 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12882 3752 3751 3682 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12881 8144 8064 3752 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12880 4410 4491 4666 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12879 8144 6867 4491 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12878 4411 4492 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12877 4666 6867 4411 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12876 8144 4901 4410 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12875 974 1024 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12874 972 1026 1019 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12873 8144 1043 972 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12872 1026 1025 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12871 8144 3708 1025 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12870 8144 1038 1024 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12869 1022 1026 974 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12868 973 1025 1022 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12867 8144 1020 973 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12866 1020 1022 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12865 1019 1025 1020 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12864 8144 1019 1043 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12863 1043 1019 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12862 3694 3832 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12861 3692 3835 3828 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12860 8144 4270 3692 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12859 3835 3836 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12858 8144 3834 3836 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12857 8144 4271 3832 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12856 3831 3835 3694 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12855 3693 3836 3831 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12854 8144 3829 3693 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12853 3829 3831 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12852 3828 3836 3829 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12851 8144 3828 4270 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12850 4270 3828 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12849 7340 8086 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12848 7340 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12847 8144 7352 7340 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12846 5507 7405 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12845 8144 7633 5507 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12844 1353 2492 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12843 7895 7966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12842 7963 7962 7895 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12841 8144 7960 7963 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12840 1470 1943 1414 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12839 8144 2616 1414 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12838 1414 2154 1470 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12837 1732 1470 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12836 3118 3570 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12835 8144 2845 3118 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12834 1547 1356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12833 8144 1553 1547 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12832 1546 957 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12831 8144 4540 1546 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12830 1545 5169 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12829 8144 1543 1545 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12828 5629 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12827 8144 7352 5629 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12826 945 942 944 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12825 944 943 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12824 8144 1119 945 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12823 1120 945 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12822 8144 6327 6563 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12821 6327 6325 6326 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12820 6324 6328 6327 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12819 8144 6325 6328 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12818 6326 6329 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12817 8144 6567 6324 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12816 6563 6327 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12815 5026 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12814 8144 5025 5026 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12813 5030 5242 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12812 8144 5872 5030 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12811 1028 5377 975 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12810 975 4651 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12809 8144 3968 1028 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12808 4658 1028 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12807 7775 7788 7776 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12806 7776 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12805 8144 8000 7775 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12804 7774 7775 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12803 2382 2847 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12802 8144 3229 2382 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12801 5885 6040 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12800 5882 6011 6038 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12799 8144 6273 5882 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12798 6011 6041 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12797 8144 8063 6041 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12796 8144 6043 6040 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12795 6010 6011 5885 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12794 5883 6041 6010 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12793 8144 6008 5883 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12792 6008 6010 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12791 6038 6041 6008 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12790 8144 6038 6273 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12789 6273 6038 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12788 7022 7033 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12787 8144 7252 7022 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12786 7517 7022 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12785 8144 6336 6334 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12784 6336 6359 6338 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12783 6337 6339 6336 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12782 8144 6359 6339 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12781 6338 7863 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12780 8144 6335 6337 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12779 6334 6336 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12778 7791 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12777 8144 5168 7791 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12776 2889 1365 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12775 8144 1550 2889 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12774 2712 2232 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12773 8144 2233 2712 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12772 7016 7025 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12771 8144 7343 7016 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12770 7329 7016 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12769 8144 7957 7746 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12768 7745 7746 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12767 8144 7979 7745 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12766 7744 7745 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12765 8144 7745 7744 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12764 7250 8000 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12763 7250 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12762 8144 7352 7250 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12761 7948 8154 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12760 7946 8157 8148 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12759 8144 8147 7946 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12758 8157 8158 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12757 8144 8166 8158 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12756 8144 8153 8154 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12755 8152 8157 7948 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12754 7947 8158 8152 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12753 8144 8150 7947 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12752 8150 8152 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12751 8148 8158 8150 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12750 8144 8148 8147 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12749 8147 8148 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12748 4083 4125 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12747 4081 4127 4120 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12746 8144 7752 4081 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12745 4127 4128 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12744 8144 8063 4128 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12743 8144 7492 4125 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12742 4124 4127 4083 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12741 4082 4128 4124 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12740 8144 4122 4082 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12739 4122 4124 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12738 4120 4128 4122 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12737 8144 4120 7752 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12736 7752 4120 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12735 5386 5388 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12734 8144 7343 5386 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12733 5553 5386 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12732 617 1798 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12731 947 7548 617 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12730 8144 6363 947 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12729 8144 4776 5232 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12728 4776 7871 4609 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12727 4608 4777 4776 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12726 8144 7871 4777 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12725 4609 7405 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12724 8144 5227 4608 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12723 5232 4776 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12722 8144 4771 4769 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12721 4771 7871 4607 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12720 4606 4773 4771 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12719 8144 7871 4773 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12718 4607 5241 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12717 8144 4770 4606 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12716 4769 4771 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12715 4602 4997 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12714 4749 5668 4602 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12713 8144 4998 4749 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12712 7627 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12711 7627 7643 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12710 8144 7888 7627 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12709 8144 7883 7627 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12708 6132 6161 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12707 6132 6133 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12706 8144 6138 6132 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12705 8144 7887 6132 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12704 5383 5606 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12703 5383 5453 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12702 8144 5938 5383 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12701 3079 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12700 3078 5907 3079 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12699 8144 6520 3078 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12698 8144 7074 7403 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12697 7074 7867 6933 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12696 6932 7077 7074 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12695 8144 7867 7077 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12694 6933 7073 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12693 8144 7270 6932 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12692 7403 7074 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12691 8144 7584 7881 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12690 7584 7867 7442 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12689 7441 7588 7584 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12688 8144 7867 7588 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12687 7442 7585 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12686 8144 7845 7441 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12685 7881 7584 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12684 5509 5740 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12683 5509 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12682 8144 6920 5509 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12681 3097 3586 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12680 3097 3735 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12679 8144 3730 3097 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12678 8144 3581 3097 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12677 8144 5558 5559 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12676 5919 6524 5528 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12675 5528 5558 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12674 5528 5559 5919 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12673 8144 5555 5528 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12672 5555 6524 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12671 5937 5940 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12670 5937 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12669 8144 6293 5937 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12668 8144 7314 5937 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12667 1856 4067 1855 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12666 3797 6796 1856 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12665 1856 2210 3797 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12664 1855 1992 1856 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12663 1855 4293 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12662 8144 2469 1855 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12661 8144 7376 7892 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12660 7376 7867 7281 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12659 7279 7282 7376 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12658 8144 7867 7282 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12657 7281 7280 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12656 8144 7581 7279 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12655 7892 7376 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12654 4312 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12653 4312 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12652 8144 6543 4312 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12651 8144 5648 4312 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12650 8144 7017 7009 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12649 7009 7006 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12648 8144 7007 7009 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12647 7321 7009 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12646 6263 6262 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12645 6261 6265 6263 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12644 8144 6260 6261 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12643 5244 5249 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12642 8144 5245 5244 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12641 5242 5244 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12640 6656 8179 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12639 8144 6654 6656 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12638 6655 6656 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12637 5179 5445 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12636 8144 6883 5179 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12635 5176 5179 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12634 7711 7955 7786 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12633 7710 7787 7711 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12632 7709 8048 7710 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12631 8144 8045 7709 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12630 8025 7786 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12629 2481 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12628 2481 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12627 8144 5447 2481 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12626 8144 4075 2481 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12625 2473 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12624 2473 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12623 8144 5648 2473 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12622 8144 5447 2473 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12621 4590 6821 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12620 4688 5406 4590 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12619 8144 6809 4688 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12618 6422 8187 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12617 6670 7408 6422 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12616 8144 7891 6670 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12615 8144 4924 4928 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12614 4925 5118 4926 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12613 4926 4924 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12612 4926 4928 4925 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12611 8144 4923 4926 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12610 4923 5118 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12609 1787 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12608 8144 7026 1787 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12607 1992 1787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12606 1302 1743 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12605 1301 1744 1302 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12604 8144 1962 1301 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12603 7799 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12602 7796 7798 7799 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12601 8144 7863 7796 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12600 8144 5390 5393 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12599 5391 7020 5392 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12598 5392 5390 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12597 5392 5393 5391 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12596 8144 5389 5392 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12595 5389 7020 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12594 2934 5496 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12593 8144 4790 2934 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12592 2932 2934 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12591 2704 2922 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12590 8144 3857 2704 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12589 2703 2704 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12588 8144 2203 1350 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12587 1350 5148 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12586 8144 1986 1350 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12585 1355 1350 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12584 8144 6293 5676 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12583 5676 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12582 5676 5940 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12581 8144 7314 5676 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12580 6138 5676 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12579 8144 7884 6174 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12578 6174 7398 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12577 6174 6893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12576 8144 7891 6174 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12575 6176 6174 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12574 8144 5942 5448 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12573 5448 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12572 5448 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12571 8144 6358 5448 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12570 5445 5448 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12569 8144 6311 4063 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12568 4063 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12567 8144 6293 4063 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12566 4061 4063 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12565 8144 2719 1387 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12564 1387 2718 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12563 8144 3857 1387 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12562 1615 1387 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12561 8144 6900 5965 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12560 5965 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12559 5965 7408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12558 8144 7891 5965 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12557 5867 5965 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12556 8144 3744 2278 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12555 2278 2334 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12554 2591 2344 2278 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12553 2277 3737 2591 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12552 2278 2589 2277 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12551 4981 4984 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12550 4977 4985 4978 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12549 8144 7867 4977 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12548 4985 4986 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12547 8144 5864 4986 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12546 8144 4983 4984 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12545 4982 4985 4981 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12544 4980 4986 4982 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12543 8144 4979 4980 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12542 4979 4982 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12541 4978 4986 4979 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12540 8144 4978 7867 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12539 7867 4978 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12538 8144 6311 1170 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12537 1170 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12536 1170 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12535 8144 4067 1170 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12534 1169 1170 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12533 8144 6900 5497 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12532 5497 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12531 5497 6893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12530 8144 7883 5497 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12529 5496 5497 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12528 8144 5447 5446 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12527 5446 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12526 8144 7353 5446 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12525 5916 5446 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12524 2454 5147 2314 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12523 2313 2698 2454 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12522 8144 4517 2313 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12521 2314 2926 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12520 7966 7965 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12519 8144 8064 7966 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12518 2175 2174 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12517 2371 4183 2175 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12516 8144 2365 2371 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12515 3115 3114 3116 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12514 3116 3552 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12513 8144 3553 3115 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12512 3112 3115 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12511 2731 2733 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12510 2727 2734 2728 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12509 8144 2964 2727 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12508 2734 2735 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12507 8144 3834 2735 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12506 8144 3267 2733 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12505 2732 2734 2731 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12504 2730 2735 2732 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12503 8144 2729 2730 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12502 2729 2732 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12501 2728 2735 2729 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12500 8144 2728 2964 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12499 2964 2728 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12498 6875 6877 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12497 6871 6879 6872 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12496 8144 6870 6871 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12495 6879 6878 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12494 8144 8166 6878 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12493 8144 6882 6877 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12492 6876 6879 6875 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12491 6874 6878 6876 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12490 8144 6873 6874 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12489 6873 6876 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12488 6872 6878 6873 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12487 8144 6872 6870 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12486 6870 6872 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12485 1791 1890 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12484 1790 1795 1791 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12483 8144 3150 1790 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12482 8144 6076 5986 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12481 5987 6801 6071 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12480 5985 6349 5987 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12479 5986 6549 5985 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12478 8144 6541 5989 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12477 5990 6520 6070 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12476 5988 6292 5990 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12475 5989 6792 5988 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12474 513 1115 516 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12473 516 1114 515 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12472 515 514 516 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12471 513 512 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12470 8144 1110 513 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12469 516 517 513 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12468 1761 515 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12467 8144 3819 3615 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12466 3615 6143 3614 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12465 3613 3614 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12464 4727 6341 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12463 4727 4728 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12462 8144 4725 4727 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12461 4744 4742 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12460 4744 5467 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12459 8144 7352 4744 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12458 6415 8179 6416 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12457 6416 7302 6415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12456 8144 6418 6416 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12455 4136 5633 4099 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12454 4099 4134 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12453 8144 4418 4136 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12452 4133 4136 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12451 4108 5003 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12450 6284 4228 4108 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12449 8144 5908 6284 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12448 3273 3275 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12447 8144 4644 3273 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12446 3751 3273 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12445 1341 1343 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12444 1337 1344 1338 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12443 8144 5443 1337 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12442 1344 1345 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12441 8144 1772 1345 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12440 8144 1526 1343 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12439 1342 1344 1341 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12438 1340 1345 1342 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12437 8144 1339 1340 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12436 1339 1342 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12435 1338 1345 1339 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12434 8144 1338 5443 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12433 5443 1338 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12432 583 652 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12431 581 651 647 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12430 8144 6520 581 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12429 651 653 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12428 8144 3708 653 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12427 8144 654 652 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12426 648 651 583 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12425 582 653 648 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12424 8144 649 582 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12423 649 648 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12422 647 653 649 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12421 8144 647 6520 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12420 6520 647 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12419 4788 4786 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12418 4788 6417 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12417 8144 4795 4788 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12416 1332 1123 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12415 8144 5641 1332 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12414 2695 1148 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12413 8144 3608 2695 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12412 2904 3378 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12411 8144 3373 2904 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12410 983 1060 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12409 981 1061 1055 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12408 8144 5394 981 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12407 1061 1062 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12406 8144 1951 1062 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12405 8144 1307 1060 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12404 1058 1061 983 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12403 982 1062 1058 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12402 8144 1056 982 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12401 1056 1058 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12400 1055 1062 1056 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12399 8144 1055 5394 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12398 5394 1055 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12397 7341 7342 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12396 8144 7343 7341 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12395 7334 7341 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12394 6538 6536 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12393 8144 6540 6538 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12392 6535 6538 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12391 2216 2924 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12390 2216 2217 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12389 8144 6359 2216 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12388 2217 2690 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12387 2217 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12386 8144 4574 2217 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12385 1889 1559 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12384 1889 1553 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12383 8144 4540 1889 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12382 1361 2262 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12381 1361 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12380 8144 4302 1361 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12379 6105 7352 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_12378 6108 6823 5921 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12377 5921 6102 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12376 8144 6100 5925 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12375 5925 6103 5924 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12374 5924 6105 6108 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12373 6108 7352 5926 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12372 5926 7528 5925 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12371 8144 6102 6100 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_12370 6829 6108 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12369 8172 7882 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12368 8172 8179 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12367 8144 7880 8172 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12366 7889 8184 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12365 7889 7888 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12364 8144 8187 7889 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12363 2722 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12362 2722 2703 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12361 8144 2894 2722 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12360 3150 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12359 3150 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12358 8144 4574 3150 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12357 4471 4583 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12356 4472 5038 4471 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12355 8144 4582 4472 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12354 3573 3763 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12353 8144 4424 3573 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12352 3571 3573 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12351 7541 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12350 7541 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12349 8144 6797 7541 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12348 8144 6549 7541 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12347 1007 1133 1134 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12346 1008 5176 1007 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12345 8144 1145 1008 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12344 1132 1134 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12343 7053 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12342 7053 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12341 8144 7354 7053 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12340 8144 8086 7053 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12339 5038 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12338 5038 6652 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12337 8144 6636 5038 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12336 8144 6921 5038 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12335 4579 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12334 4579 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12333 8144 4575 4579 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12332 8144 4302 4579 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12331 5037 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12330 5037 6636 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12329 8144 6396 5037 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12328 8144 6921 5037 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12327 3759 8139 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12326 3759 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12325 8144 4172 3759 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12324 8144 7749 7496 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12323 7496 7518 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12322 7496 7725 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12321 8144 7724 7496 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12320 7730 7496 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12319 5014 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12318 8144 6396 5014 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12317 5013 5014 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12316 7048 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12315 7048 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12314 8144 7354 7048 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12313 8144 8071 7048 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12312 1587 5148 1434 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12311 1433 2698 1587 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12310 8144 4518 1433 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12309 1434 2926 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_12308 1866 1892 2025 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12307 1867 1893 1866 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12306 8144 2700 1867 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12305 2942 2025 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12304 2843 3759 2756 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12303 2756 4166 2843 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12302 8144 4510 2756 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12301 3675 3720 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12300 3722 4492 3675 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12299 8144 8064 3722 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12298 6056 6489 5980 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12297 8144 6055 5980 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12296 5980 6480 6056 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12295 6786 6056 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12294 3358 3610 3215 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12293 3215 4556 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12292 8144 3788 3358 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12291 3356 3358 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12290 8144 786 785 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12289 4068 785 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12288 8144 785 4068 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12287 8144 785 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12286 8144 785 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12285 8144 786 787 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12284 4573 787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12283 8144 787 4573 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12282 8144 787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12281 8144 787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12280 8144 576 577 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12279 786 577 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12278 8144 577 786 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12277 8144 577 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12276 8144 577 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12275 8144 3179 2489 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12274 6543 2489 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12273 8144 2489 6543 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12272 8144 2489 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12271 8144 2489 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12270 8144 3179 2726 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12269 6797 2726 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12268 8144 2726 6797 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12267 8144 2726 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12266 8144 2726 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12265 8144 3179 2720 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12264 7356 2720 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12263 8144 2720 7356 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12262 8144 2720 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12261 8144 2720 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12260 8144 3179 3180 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12259 4051 3180 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12258 8144 3180 4051 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12257 8144 3180 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12256 8144 3180 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12255 8144 2490 2491 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12254 3179 2491 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12253 8144 2491 3179 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12252 8144 2491 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12251 8144 2491 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12250 552 3622 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12249 8144 1150 552 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12248 551 552 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12247 1318 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12246 8144 1317 1318 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12245 1956 1318 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12244 8144 6658 6411 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12243 6411 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12242 8144 7130 6411 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12241 6410 6411 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12240 2716 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12239 8144 7051 2716 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12238 2938 2716 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12237 6518 6835 6435 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12236 6435 7073 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12235 8144 6794 6518 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12234 6517 6518 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12233 8144 5483 5484 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12232 5484 5654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12231 5484 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12230 8144 7500 5484 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12229 7880 5484 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12228 3420 3415 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12227 8144 4311 3420 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12226 3416 3420 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12225 8144 6802 2449 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12224 2449 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12223 8144 2687 2449 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12222 2696 2449 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12221 8144 4208 4210 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12220 4210 4212 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12219 8144 4206 4210 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12218 4207 4210 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12217 5945 6131 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12216 5941 6025 6125 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12215 8144 6127 5941 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12214 6025 6130 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12213 8144 7821 6130 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12212 8144 6128 6131 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12211 6024 6025 5945 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12210 5943 6130 6024 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12209 8144 6022 5943 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12208 6022 6024 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12207 6125 6130 6022 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12206 8144 6125 6127 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12205 6127 6125 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12204 8144 5624 1162 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12203 1162 1565 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12202 1162 5483 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12201 8144 3857 1162 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12200 1381 1162 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12199 2687 1799 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12198 2690 5940 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12197 774 2964 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12196 7581 7845 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12195 7270 7572 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12194 7076 7272 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12193 8144 7619 7618 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12192 7618 8186 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12191 8144 7869 7618 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12190 7887 7618 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12189 8144 5147 3346 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12188 3346 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12187 3346 7343 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12186 8144 5148 3346 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12185 3794 3346 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12184 8144 7026 4027 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12183 4027 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12182 4027 4572 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12181 8144 5003 4027 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12180 6090 4027 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12179 4155 4143 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12178 8144 3986 4155 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12177 881 882 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12176 876 883 877 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12175 8144 1304 876 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12174 883 884 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12173 8144 1951 884 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12172 8144 885 882 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12171 880 883 881 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12170 878 884 880 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12169 8144 879 878 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12168 879 880 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12167 877 884 879 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12166 8144 877 1304 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12165 1304 877 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12164 7370 7778 7269 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12163 7269 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12162 8144 7863 7370 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12161 7367 7370 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12160 5653 6883 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12159 4134 5563 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12158 2789 5387 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12157 5380 5394 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12156 8144 2492 236 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12155 236 1799 369 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12154 8144 2964 580 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12153 580 2968 579 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12152 8144 2471 2033 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12151 2033 1902 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12150 2033 1899 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12149 8144 2035 2033 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12148 3642 2033 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12147 3546 3316 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12146 8144 3229 3546 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12145 7951 8168 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12144 7949 8167 8161 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12143 8144 8159 7949 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12142 8167 8170 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12141 8144 8166 8170 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12140 8144 8173 8168 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12139 8165 8167 7951 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12138 7950 8170 8165 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12137 8144 8162 7950 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12136 8162 8165 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12135 8161 8170 8162 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12134 8144 8161 8159 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12133 8159 8161 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12132 7043 8071 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12131 7043 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12130 8144 7041 7043 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12129 5156 6294 5057 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12128 5057 7056 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12127 8144 5162 5156 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12126 5416 5156 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12125 8144 2906 1861 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12124 1861 2011 2004 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12123 2005 2004 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12122 8144 2906 1860 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12121 1860 2006 2002 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_12120 2003 2002 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12119 1346 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12118 8144 1335 1346 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12117 7245 7955 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12116 7729 7747 7245 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12115 8144 7319 7729 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12114 3327 3763 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12113 8144 4424 3327 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12112 6771 6773 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12111 6767 6774 6768 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12110 8144 6775 6767 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12109 6774 6776 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12108 8144 8063 6776 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12107 8144 6780 6773 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12106 6772 6774 6771 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12105 6769 6776 6772 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12104 8144 6770 6769 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12103 6770 6772 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12102 6768 6776 6770 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12101 8144 6768 6775 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12100 6775 6768 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12099 8144 6094 6319 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12098 6094 6095 5994 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12097 5993 6097 6094 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12096 8144 6095 6097 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12095 5994 6096 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12094 8144 6344 5993 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12093 6319 6094 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12092 8144 5918 6096 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12091 5918 5842 5843 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12090 5841 5844 5918 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12089 8144 5842 5844 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12088 5843 7549 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12087 8144 6292 5841 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12086 6096 5918 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12085 5053 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12084 5132 5907 5053 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12083 8144 6076 5132 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12082 2924 2469 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12081 8144 7051 2924 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12080 1306 5828 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12079 8144 1313 1306 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12078 2213 2682 2211 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12077 2211 2210 2212 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12076 2212 7051 2213 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12075 2213 2894 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12074 8144 4067 2213 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12073 2679 2212 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12072 2648 4947 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12071 8144 3134 2648 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12070 7943 8133 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12069 7941 8134 8127 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12068 8144 8125 7941 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12067 8134 8135 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12066 8144 8166 8135 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12065 8144 8130 8133 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12064 8132 8134 7943 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12063 7942 8135 8132 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12062 8144 8128 7942 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12061 8128 8132 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12060 8127 8135 8128 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12059 8144 8127 8125 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12058 8125 8127 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12057 6058 6784 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12056 8144 6785 6058 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12055 6503 6058 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12054 5407 5414 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12053 8144 5616 5407 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12052 6785 5407 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12051 6548 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12050 8144 7352 6548 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12049 7760 6548 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12048 8144 6356 6581 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12047 6356 6362 6355 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12046 6354 6357 6356 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12045 8144 6362 6357 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12044 6355 6576 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12043 8144 6353 6354 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12042 6581 6356 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12041 8144 6119 6353 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12040 6119 6359 5998 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12039 5997 6120 6119 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12038 8144 6359 6120 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12037 5998 7777 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12036 8144 6347 5997 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_12035 6353 6119 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12034 1996 2469 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12033 8144 4306 1996 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12032 7877 7891 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12031 7877 7643 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12030 8144 7888 7877 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12029 7017 8021 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12028 7017 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12027 8144 7352 7017 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12026 2798 2796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12025 2798 3586 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12024 8144 3581 2798 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12023 8144 3542 2798 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12022 3143 3146 3142 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12021 3142 4007 3143 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12020 8144 4510 3142 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12019 1834 1918 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12018 1832 1917 1913 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12017 8144 5906 1832 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12016 1917 1919 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12015 8144 3708 1919 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_12014 8144 3508 1918 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12013 1878 1917 1834 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12012 1833 1919 1878 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12011 8144 1877 1833 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12010 1877 1878 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12009 1913 1919 1877 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_12008 8144 1913 5906 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12007 5906 1913 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_12006 7312 7313 7242 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12005 7242 7518 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12004 8144 7314 7312 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12003 7486 7312 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_12002 4651 5606 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12001 4651 5384 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_12000 8144 6792 4651 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11999 8144 5888 5551 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11998 8144 7500 5552 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11997 5551 5552 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11996 3393 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11995 3393 5654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11994 8144 5483 3393 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11993 8144 4461 3393 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11992 8144 4173 2615 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11991 2615 4172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11990 8144 7585 2615 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11989 2614 2615 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11988 8144 4022 4023 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11987 6152 4023 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11986 8144 4023 6152 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11985 8144 4023 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11984 8144 4023 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11983 8144 3792 3793 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11982 5961 3793 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11981 8144 3793 5961 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11980 8144 3793 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11979 8144 3793 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11978 8144 6152 6153 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11977 8166 6153 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11976 8144 6153 8166 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11975 8144 6153 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11974 8144 6153 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11973 8144 6152 6151 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11972 7821 6151 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11971 8144 6151 7821 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11970 8144 6151 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11969 8144 6151 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11968 8144 6152 5963 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11967 5864 5963 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11966 8144 5963 5864 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11965 8144 5963 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11964 8144 5963 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11963 8144 5961 5962 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11962 5863 5962 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11961 8144 5962 5863 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11960 8144 5962 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11959 8144 5962 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11958 8144 6152 6069 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11957 8063 6069 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11956 8144 6069 8063 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11955 8144 6069 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11954 8144 6069 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11953 8144 6152 6068 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11952 6067 6068 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11951 8144 6068 6067 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11950 8144 6068 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11949 8144 6068 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11948 8144 1446 1447 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11947 5558 5453 1411 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11946 1411 1446 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11945 1411 1447 5558 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11944 8144 1443 1411 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11943 1443 5453 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11942 8178 8182 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11941 8144 8175 8178 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11940 8176 8178 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11939 8144 4955 4232 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11938 4233 4232 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11937 8144 4230 4233 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11936 4530 4233 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11935 8144 4233 4530 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11934 8144 2968 792 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11933 789 792 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11932 8144 2964 789 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11931 791 789 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11930 8144 789 791 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11929 3073 2957 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11928 3073 3860 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11927 8144 2958 3073 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11926 3622 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11925 3622 5654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11924 8144 5483 3622 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11923 8144 5015 3622 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11922 8144 3293 2613 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11921 2613 3566 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11920 8144 3744 2613 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11919 2612 2613 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11918 3730 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11917 3730 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11916 8144 4167 3730 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11915 8144 6273 3730 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11914 8144 5603 5909 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11913 8144 7314 5605 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11912 5909 5605 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11911 5706 5868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11910 5706 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11909 8144 6632 5706 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11908 8144 7130 5706 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11907 6458 6629 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11906 6617 6615 6458 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11905 8144 6614 6617 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11904 4649 5379 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11903 8144 4647 4649 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11902 4648 4649 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11901 4935 5429 4938 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11900 4936 7787 4935 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11899 4937 8048 4936 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11898 8144 8045 4937 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11897 4934 4938 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11896 8144 3787 3621 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11895 3639 5453 3620 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11894 3620 3787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11893 3620 3621 3639 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11892 8144 3619 3620 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11891 3619 5453 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11890 8144 4921 4922 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11889 4924 7056 4920 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11888 4920 4921 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11887 4920 4922 4924 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11886 8144 4919 4920 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11885 4919 7056 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11884 7433 7559 7432 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11883 7432 7548 7552 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11882 7552 7550 7433 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11881 7433 7804 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11880 8144 7554 7433 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11879 7547 7552 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11878 5138 5140 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11877 8144 5408 5138 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11876 5136 5138 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11875 3609 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11874 8144 5168 3609 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11873 3801 3609 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11872 1781 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11871 8144 5147 1781 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11870 1780 1781 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11869 575 2964 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11868 8144 2968 575 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11867 574 575 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11866 2459 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11865 8144 2718 2459 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11864 2706 2459 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11863 5984 6267 5983 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11862 6301 8008 5984 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11861 5984 6285 6301 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11860 5983 6286 5984 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11859 5983 6520 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11858 8144 6284 5983 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11857 3306 3993 3203 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11856 3203 3987 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11855 8144 3315 3306 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11854 3303 3306 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11853 4005 5406 4006 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11852 4006 7056 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11851 8144 6812 4005 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11850 4003 4005 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11849 8144 2886 2411 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11848 2411 2413 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11847 8144 2407 2411 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11846 2408 2411 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11845 6844 6846 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11844 6839 6848 6840 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11843 8144 6838 6839 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11842 6848 6847 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11841 8144 7821 6847 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11840 8144 6843 6846 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11839 6845 6848 6844 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11838 6842 6847 6845 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11837 8144 6841 6842 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11836 6841 6845 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11835 6840 6847 6841 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11834 8144 6840 6838 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11833 6838 6840 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11832 6888 6890 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11831 6884 6892 6885 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11830 8144 6883 6884 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11829 6892 6891 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11828 8144 8166 6891 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11827 8144 6899 6890 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11826 6889 6892 6888 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11825 6887 6891 6889 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11824 8144 6886 6887 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11823 6886 6889 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11822 6885 6891 6886 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11821 8144 6885 6883 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11820 6883 6885 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11819 4597 4722 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11818 4721 7352 4597 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11817 8144 4739 4721 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11816 8144 8187 5493 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11815 5493 6900 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11814 8144 7883 5493 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11813 5492 5493 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11812 7407 7408 7306 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11811 7306 7881 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11810 8144 7891 7407 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11809 7305 7407 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11808 3133 3582 3066 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11807 8144 3579 3066 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11806 3066 3356 3133 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11805 3552 3133 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11804 2171 2170 2173 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11803 2173 4189 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11802 8144 2375 2171 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11801 2168 2171 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11800 590 669 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11799 588 668 664 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11798 8144 677 588 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11797 668 670 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11796 8144 1951 670 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11795 8144 671 669 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11794 665 668 590 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11793 589 670 665 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11792 8144 666 589 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11791 666 665 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11790 664 670 666 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11789 8144 664 677 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11788 677 664 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11787 7770 7774 8006 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11786 7769 7767 7770 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11785 8144 7768 7769 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11784 1002 1743 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11783 1052 1744 1002 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11782 8144 8045 1052 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11781 8144 4295 1605 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11780 1605 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11779 1605 4293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11778 8144 5648 1605 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11777 1897 1605 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11776 4802 5737 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11775 8144 5740 4802 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11774 7728 7738 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11773 8144 7730 7728 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11772 8144 5453 2318 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11771 8144 7314 1282 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11770 2318 1282 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11769 6392 6393 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11768 6387 6395 6388 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11767 8144 6398 6387 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11766 6395 6394 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11765 8144 8166 6394 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11764 8144 6401 6393 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11763 6390 6395 6392 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11762 6389 6394 6390 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11761 8144 6391 6389 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11760 6391 6390 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11759 6388 6394 6391 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11758 8144 6388 6398 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11757 6398 6388 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11756 6665 7408 6465 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11755 6465 7884 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11754 8144 7891 6665 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11753 6914 6665 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11752 1846 2179 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11751 2172 2178 1846 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11750 8144 3148 2172 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11749 3556 3780 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11748 8144 4255 3556 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11747 2827 3348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11746 2827 3989 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11745 8144 3990 2827 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11744 2187 2190 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11743 2183 2191 2184 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11742 8144 5143 2183 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11741 2191 2192 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11740 8144 3708 2192 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11739 8144 2189 2190 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11738 2188 2191 2187 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11737 2186 2192 2188 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11736 8144 2185 2186 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11735 2185 2188 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11734 2184 2192 2185 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11733 8144 2184 5143 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11732 5143 2184 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11731 903 1123 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11730 8144 1115 903 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11729 3629 3624 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11728 8144 3253 3629 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11727 7743 7754 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11726 8144 7742 7743 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11725 3989 7349 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11724 3989 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11723 8144 4172 3989 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11722 3089 3088 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11721 3080 3083 3081 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11720 8144 6792 3080 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11719 3083 3091 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11718 8144 3708 3091 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11717 8144 3962 3088 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11716 3085 3083 3089 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11715 3086 3091 3085 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11714 8144 3084 3086 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11713 3084 3085 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11712 3081 3091 3084 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11711 8144 3081 6792 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11710 6792 3081 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11709 6299 6298 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11708 8144 7343 6299 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11707 6297 6299 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11706 5502 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11705 5502 5971 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11704 8144 6909 5502 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11703 939 1123 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11702 8144 1114 939 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11701 2693 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11700 2693 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11699 8144 4068 2693 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11698 5238 6652 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11697 8144 6172 5238 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11696 1733 3958 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11695 1735 2672 1731 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11694 1731 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11693 8144 1730 1737 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11692 1737 1732 1734 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11691 1734 1733 1735 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11690 1735 3958 1736 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11689 1736 2155 1737 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11688 8144 3556 1730 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11687 1729 1735 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11686 1938 3958 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11685 1941 3009 1840 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11684 1840 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11683 8144 1935 1843 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11682 1843 1936 1841 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11681 1841 1938 1941 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11680 1941 3958 1842 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11679 1842 2154 1843 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11678 8144 3556 1935 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11677 2132 1941 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11676 3105 3989 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11675 8144 3990 3105 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11674 3104 3105 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11673 1407 1515 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11672 1405 1517 1510 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11671 8144 5419 1405 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11670 1517 1518 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11669 8144 1772 1518 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11668 8144 1519 1515 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11667 1514 1517 1407 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11666 1406 1518 1514 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11665 8144 1512 1406 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11664 1512 1514 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11663 1510 1518 1512 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11662 8144 1510 5419 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11661 5419 1510 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11660 7318 6472 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11659 7318 6477 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11658 8144 6478 7318 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11657 8144 6473 7318 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11656 3076 6473 3075 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11655 3075 6472 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11654 8144 8064 3076 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11653 6087 3076 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11652 5724 7130 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11651 5724 6176 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11650 8144 6921 5724 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11649 8144 7835 7264 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11648 8144 7957 7265 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11647 7264 7265 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11646 4582 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11645 4582 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11644 8144 4575 4582 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11643 8144 4306 4582 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11642 6463 7398 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11641 6652 7884 6463 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11640 8144 7891 6652 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11639 1319 1965 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11638 1752 1964 1319 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11637 8144 3148 1752 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11636 8144 4173 2014 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11635 2014 4172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11634 8144 7549 2014 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11633 2156 2014 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11632 1714 2144 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11631 1715 3958 1713 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11630 1713 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11629 8144 1712 1717 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11628 1717 1925 1716 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11627 1716 1714 1715 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11626 1715 2144 1718 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11625 1718 2605 1717 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11624 8144 3556 1712 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11623 1711 1715 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11622 1461 2144 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11621 1463 1467 1395 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11620 1395 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11619 8144 1459 1398 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11618 1398 1932 1396 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11617 1396 1461 1463 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11616 1463 2144 1397 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11615 1397 2608 1398 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11614 8144 3556 1459 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_11613 2136 1463 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11612 7342 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11611 7342 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11610 8144 7354 7342 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11609 8144 7824 7342 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11608 2927 2924 2778 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11607 2778 2926 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11606 8144 2925 2927 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11605 3405 2927 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11604 8144 7250 7005 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11603 7005 7002 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11602 8144 7011 7005 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11601 7508 7005 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11600 8144 1796 1797 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11599 1797 1891 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11598 8144 6363 1797 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11597 4236 1797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11596 1698 2698 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11595 1805 2924 1698 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11594 1697 1806 1805 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11593 8144 2926 1697 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11592 2232 1805 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11591 3220 3251 3392 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11590 3221 3252 3220 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11589 8144 3250 3221 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11588 3409 3392 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11587 5839 6090 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11586 5838 6089 5839 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11585 8144 6344 5838 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11584 8144 3100 3093 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11583 3720 3095 3096 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11582 3096 3100 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11581 3096 3093 3720 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11580 8144 3094 3096 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11579 3094 3095 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11578 8144 4076 3855 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11577 7026 3855 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11576 8144 3855 7026 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11575 8144 3855 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11574 8144 3855 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11573 8144 4076 4077 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11572 6609 4077 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11571 8144 4077 6609 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11570 8144 4077 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11569 8144 4077 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11568 8144 4076 4065 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11567 7354 4065 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11566 8144 4065 7354 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11565 8144 4065 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11564 8144 4065 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11563 8144 3662 3663 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11562 4076 3663 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11561 8144 3663 4076 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11560 8144 3663 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11559 8144 3663 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11558 8144 568 567 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11557 4293 567 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11556 8144 567 4293 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11555 8144 567 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11554 8144 567 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11553 8144 568 569 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11552 4302 569 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11551 8144 569 4302 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11550 8144 569 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11549 8144 569 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11548 8144 568 566 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11547 4572 566 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11546 8144 566 4572 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11545 8144 566 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11544 8144 566 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11543 8144 375 376 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11542 568 376 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11541 8144 376 568 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11540 8144 376 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11539 8144 376 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11538 5537 5653 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11537 5922 5641 5537 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11536 8144 5642 5922 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11535 5716 5870 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11534 8144 5728 5716 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11533 5967 5716 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11532 8144 7398 6910 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11531 6910 7884 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11530 8144 7883 6910 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11529 6909 6910 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11528 7427 7750 7532 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11527 7426 7787 7427 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11526 7425 8048 7426 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11525 8144 8045 7425 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11524 7566 7532 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11523 4435 6304 4515 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11522 4436 7787 4435 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11521 4434 8048 4436 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11520 8144 8045 4434 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11519 4433 4515 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11518 7736 7962 7735 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11517 7735 7734 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11516 8144 7957 7736 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11515 7733 7736 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11514 8144 782 571 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11513 4306 571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11512 8144 571 4306 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11511 8144 571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11510 8144 571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11509 8144 782 570 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11508 4067 570 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11507 8144 570 4067 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11506 8144 570 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11505 8144 570 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11504 8144 782 783 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11503 5624 783 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11502 8144 783 5624 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11501 8144 783 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11500 8144 783 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11499 8144 378 377 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11498 782 377 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11497 8144 377 782 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11496 8144 377 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11495 8144 377 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11494 8144 1190 1191 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11493 4574 1191 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11492 8144 1191 4574 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11491 8144 1191 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11490 8144 1191 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11489 8144 1190 971 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11488 5648 971 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11487 8144 971 5648 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11486 8144 971 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11485 8144 971 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11484 8144 1190 967 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11483 4167 967 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11482 8144 967 4167 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11481 8144 967 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11480 8144 967 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11479 8144 791 788 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11478 1190 788 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11477 8144 788 1190 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11476 8144 788 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11475 8144 788 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11474 6305 6304 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11473 6477 7747 6305 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11472 8144 6535 6477 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11471 8144 7892 6638 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11470 6638 7408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11469 8144 7883 6638 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11468 6654 6638 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11467 2231 2232 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11466 8144 2233 2231 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11465 2240 2231 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11464 2472 2469 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11463 8144 4306 2472 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11462 2943 2472 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11461 2724 2722 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11460 8144 2723 2724 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11459 3415 2724 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11458 8144 4049 3825 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11457 4295 3825 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11456 8144 3825 4295 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11455 8144 3825 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11454 8144 3825 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11453 8144 4049 4050 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11452 4575 4050 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11451 8144 4050 4575 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11450 8144 4050 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11449 8144 4050 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11448 8144 4045 4046 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11447 4049 4046 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11446 8144 4046 4049 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11445 8144 4046 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11444 8144 4046 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11443 6951 7059 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11442 7369 7058 6951 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11441 8144 7062 7369 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11440 1865 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11439 2017 2203 1865 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11438 1864 2227 2017 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11437 8144 2698 1864 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11436 2235 2017 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11435 5974 7893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11434 8144 8184 5974 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11433 5878 5974 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11432 2444 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11431 8144 4574 2444 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11430 2688 2444 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11429 8144 2719 1386 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11428 1386 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11427 8144 3857 1386 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11426 1389 1386 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11425 8144 359 347 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11424 347 1150 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11423 8144 4558 347 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11422 343 347 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11421 8144 7954 7960 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11420 8144 8064 6468 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11419 7960 6468 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11418 991 1086 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11417 989 1085 1080 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11416 8144 1758 989 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11415 1085 1087 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11414 8144 1772 1087 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11413 8144 1091 1086 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11412 1083 1085 991 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11411 990 1087 1083 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11410 8144 1081 990 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11409 1081 1083 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11408 1080 1087 1081 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11407 8144 1080 1758 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11406 1758 1080 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11405 5543 6618 5682 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11404 5542 6398 5543 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11403 8144 6141 5542 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11402 5539 6127 5665 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11401 5538 5664 5539 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11400 8144 6143 5538 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11399 4541 4749 4450 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11398 4450 4987 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11397 8144 4540 4541 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11396 4449 4541 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11395 8144 7619 6908 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11394 6908 6907 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11393 6908 8186 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11392 8144 8184 6908 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11391 6906 6908 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11390 5634 5633 5533 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11389 5533 5632 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11388 8144 7547 5634 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11387 5912 5634 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11386 5129 5419 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11385 5567 5571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11384 5632 5435 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11383 2609 2809 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11382 2608 3320 2609 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11381 8144 3315 2608 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11380 2831 3310 2754 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11379 2754 2833 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11378 8144 2830 2831 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11377 4498 2831 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11376 5861 5957 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11375 5859 5958 5952 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11374 8144 6143 5859 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11373 5958 5960 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11372 8144 7821 5960 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11371 8144 6386 5957 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11370 5955 5958 5861 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11369 5860 5960 5955 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11368 8144 5954 5860 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11367 5954 5955 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11366 5952 5960 5954 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11365 8144 5952 6143 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11364 6143 5952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11363 1794 2439 1795 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11362 1793 1792 1794 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11361 8144 2003 1793 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11360 948 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11359 8144 1372 948 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11358 5444 5443 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11357 5421 5143 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11356 7758 7979 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11355 8009 8008 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11354 7955 7954 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11353 7802 3077 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11352 8144 4293 1393 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11351 1393 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11350 1393 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11349 8144 4075 1393 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11348 1617 1393 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11347 8144 6797 2255 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11346 2255 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11345 2255 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11344 8144 5942 2255 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11343 2254 2255 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11342 3748 4511 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11341 8144 4512 3748 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11340 996 1102 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11339 994 1104 1097 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11338 8144 1335 994 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11337 1104 1105 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11336 8144 1772 1105 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11335 8144 1330 1102 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11334 1101 1104 996 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11333 995 1105 1101 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11332 8144 1099 995 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11331 1099 1101 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11330 1097 1105 1099 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11329 8144 1097 1335 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11328 1335 1097 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11327 4459 4566 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11326 4457 4567 4564 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11325 8144 4734 4457 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11324 4567 4569 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11323 8144 5864 4569 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11322 8144 4570 4566 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11321 4565 4567 4459 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11320 4458 4569 4565 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11319 8144 4568 4458 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11318 4568 4565 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11317 4564 4569 4568 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11316 8144 4564 4734 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11315 4734 4564 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11314 4529 3370 3219 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_11313 3218 5624 4529 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_11312 8144 4302 3218 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_11311 3219 3371 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_11310 4963 4537 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11309 8144 4727 4963 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11308 4766 6383 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11307 8144 4635 4766 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11306 4730 4230 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11305 3686 4021 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11304 4193 7788 3686 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11303 8144 6792 4193 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11302 8144 2129 2126 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11301 2129 6867 2130 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11300 2128 2131 2129 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11299 8144 6867 2131 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11298 2130 2133 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11297 8144 2127 2128 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11296 2126 2129 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11295 3562 4685 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11294 8144 2361 3562 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11293 7336 7824 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11292 7336 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11291 8144 7352 7336 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11290 8144 6352 6347 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11289 6352 6358 6351 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11288 6348 6350 6352 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11287 8144 6358 6350 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11286 6351 6349 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11285 8144 6586 6348 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11284 6347 6352 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11283 2935 5496 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11282 8144 4790 2935 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11281 1753 4437 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11280 8144 1752 1753 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11279 2636 2635 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11278 8144 3137 2636 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11277 1290 2595 1288 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11276 1288 1287 1289 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11275 1289 1929 1290 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11274 1290 1451 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11273 8144 2132 1290 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11272 1296 1289 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11271 6429 6497 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11270 6427 6498 6490 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11269 8144 6489 6427 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11268 6498 6499 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11267 8144 8063 6499 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11266 8144 6495 6497 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11265 6494 6498 6429 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11264 6428 6499 6494 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11263 8144 6492 6428 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11262 6492 6494 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11261 6490 6499 6492 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11260 8144 6490 6489 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11259 6489 6490 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11258 4109 4234 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11257 4537 4447 4109 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11256 8144 5449 4537 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11255 8144 6376 6374 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11254 6376 6383 6380 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11253 6377 6379 6376 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11252 8144 6383 6379 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11251 6380 6378 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11250 8144 6375 6377 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11249 6374 6376 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11248 5042 7149 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11247 5042 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11246 8144 7887 5042 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11245 4929 5600 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11244 8144 4927 4929 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11243 2199 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11242 8144 5147 2199 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11241 3788 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11240 3788 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11239 8144 7354 3788 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11238 8144 3787 3788 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11237 7938 8115 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11236 7936 8116 8110 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11235 8144 8119 7936 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11234 8116 8117 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11233 8144 8166 8117 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11232 8144 8118 8115 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11231 8113 8116 7938 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11230 7937 8117 8113 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11229 8144 8111 7937 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11228 8111 8113 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11227 8110 8117 8111 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11226 8144 8110 8119 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11225 8119 8110 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11224 7795 7794 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11223 8144 7796 7795 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11222 7793 7795 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11221 5531 5588 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11220 5589 6785 5531 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11219 8144 5587 5589 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11218 5927 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11217 5927 5854 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11216 8144 5654 5927 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11215 8144 6796 5927 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11214 8144 5481 5478 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11213 5481 7871 5480 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11212 5479 5482 5481 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11211 8144 7871 5482 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11210 5480 5712 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11209 8144 5664 5479 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11208 5478 5481 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11207 8144 4258 4254 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11206 4258 7871 4093 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11205 4092 4259 4258 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11204 8144 7871 4259 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11203 4093 5013 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11202 8144 4255 4092 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11201 4254 4258 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11200 8144 4762 4759 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11199 4762 7871 4605 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11198 4604 4764 4762 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11197 8144 7871 4764 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11196 4605 5495 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11195 8144 4760 4604 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11194 4759 4762 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11193 8144 7137 5723 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11192 5722 5723 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11191 8144 5968 5722 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11190 5720 5722 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11189 8144 5722 5720 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11188 8144 3356 3334 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11187 3334 3581 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11186 8144 3582 3334 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11185 3744 3334 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11184 8144 5199 5196 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11183 5199 7871 5065 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11182 5064 5200 5199 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11181 8144 7871 5200 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11180 5065 6154 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11179 8144 5197 5064 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11178 5196 5199 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11177 6948 7020 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11176 7782 7058 6948 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11175 8144 7025 7782 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11174 8144 1381 1383 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11173 1383 1384 1382 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11172 2249 1382 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11171 8144 1168 1014 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11170 1014 1169 1166 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11169 1589 1166 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11168 1430 1571 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11167 3171 1570 1430 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11166 8144 7550 3171 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11165 7137 7630 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11164 7137 7884 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11163 8144 7888 7137 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11162 8144 8184 7137 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11161 4476 5740 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11160 4476 5737 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11159 8144 4790 4476 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11158 4228 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11157 4228 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11156 8144 6609 4228 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11155 1863 2220 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11154 2013 2011 1863 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11153 8144 8159 2013 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11152 5979 6786 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11151 6278 6503 5979 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11150 8144 7500 6278 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11149 6360 6364 6362 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11148 8144 6363 6364 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11147 6361 6607 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11146 6362 6363 6361 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11145 8144 6359 6360 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11144 8144 6500 6046 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11143 6046 6051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11142 6046 6786 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11141 8144 6503 6046 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11140 6473 6046 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11139 8144 2875 2879 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11138 2877 2873 2761 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11137 2761 2875 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11136 2761 2879 2877 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11135 8144 2876 2761 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11134 2876 2873 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_11133 8144 7892 7641 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11132 7641 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11131 8144 7891 7641 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11130 7639 7641 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11129 2900 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11128 8144 7356 2900 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11127 2898 2900 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11126 1591 3253 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11125 8144 1590 1591 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11124 1819 1591 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11123 1010 4067 1009 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11122 1009 1353 1143 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11121 1143 1140 1010 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11120 1010 7051 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11119 8144 2894 1010 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11118 1139 1143 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11117 5131 5633 5055 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11116 5055 5129 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11115 8144 6530 5131 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11114 5151 5131 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11113 8144 7643 7636 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11112 7636 7888 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11111 8144 7891 7636 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11110 7633 7636 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11109 8144 3260 3185 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11108 3185 3858 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11107 8144 3184 3185 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11106 3192 3185 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11105 8144 4230 4028 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11104 4028 4538 4029 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11103 3204 3987 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11102 3307 3993 3204 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11101 8144 3315 3307 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11100 6813 6835 6814 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11099 6814 7612 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11098 8144 7342 6813 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11097 6812 6813 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_11096 542 545 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11095 539 546 540 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11094 8144 739 539 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11093 546 547 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11092 8144 3834 547 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11091 8144 740 545 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11090 543 546 542 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11089 544 547 543 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11088 8144 541 544 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11087 541 543 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11086 540 547 541 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11085 8144 540 739 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11084 739 540 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11083 6408 6909 6406 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11082 6409 6912 6408 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11081 6408 6407 6409 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11080 6406 7135 6408 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11079 6406 6410 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11078 8144 6647 6406 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11077 8144 7630 7132 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11076 7132 7893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11075 8144 8184 7132 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11074 7130 7132 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11073 2774 2919 3636 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11072 2773 2918 2774 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11071 8144 3251 2773 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11070 8144 1619 1613 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11069 1613 1611 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11068 8144 2448 1613 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11067 3863 1613 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11066 6858 6860 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11065 6854 6861 6855 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11064 8144 6864 6854 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11063 6861 6862 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11062 8144 7821 6862 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11061 8144 6863 6860 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11060 6859 6861 6858 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11059 6857 6862 6859 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11058 8144 6856 6857 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11057 6856 6859 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11056 6855 6862 6856 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11055 8144 6855 6864 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11054 6864 6855 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11053 4523 4704 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11052 4520 4627 4702 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11051 8144 4714 4520 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11050 4627 4706 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11049 8144 8063 4706 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11048 8144 7549 4704 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11047 4626 4627 4523 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11046 4522 4706 4626 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11045 8144 4624 4522 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11044 4624 4626 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11043 4702 4706 4624 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11042 8144 4702 4714 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11041 4714 4702 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11040 7422 7525 7772 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11039 7421 7459 7422 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11038 8144 7529 7421 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11037 86 88 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11036 82 89 83 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11035 8144 268 82 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11034 89 90 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11033 8144 1951 90 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11032 8144 91 88 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11031 87 89 86 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11030 84 90 87 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11029 8144 85 84 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11028 85 87 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11027 83 90 85 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11026 8144 83 268 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11025 268 83 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11024 5526 5688 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11023 5524 5690 5683 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11022 8144 6141 5524 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11021 5690 5691 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11020 8144 5864 5691 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_11019 8144 5704 5688 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11018 5687 5690 5526 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11017 5525 5691 5687 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11016 8144 5685 5525 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11015 5685 5687 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11014 5683 5691 5685 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_11013 8144 5683 6141 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11012 6141 5683 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11011 5530 7020 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11010 5823 6294 5530 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11009 8144 5825 5823 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11008 5923 6363 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11007 5923 6359 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11006 8144 5908 5923 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11005 8144 6145 5995 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11004 5995 6618 6111 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_11003 6112 6111 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_11002 8015 8006 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11001 8144 8004 8015 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_11000 6000 7881 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10999 6172 7408 6000 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10998 8144 7891 6172 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10997 3597 3600 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10996 3592 3601 3593 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10995 8144 3787 3592 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10994 3601 3599 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10993 8144 3834 3599 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10992 8144 3596 3600 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10991 3598 3601 3597 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10990 3594 3599 3598 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10989 8144 3595 3594 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10988 3595 3598 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10987 3593 3599 3595 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10986 8144 3593 3787 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10985 3787 3593 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10984 3528 3529 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10983 3524 3531 3523 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10982 8144 6541 3524 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10981 3531 3530 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10980 8144 3708 3530 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10979 8144 3718 3529 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10978 3526 3531 3528 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10977 3527 3530 3526 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10976 8144 3525 3527 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10975 3525 3526 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10974 3523 3530 3525 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10973 8144 3523 6541 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10972 6541 3523 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10971 7727 7724 7726 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10970 7726 7725 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10969 8144 7957 7727 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10968 7723 7727 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10967 5845 6112 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10966 6103 5919 5845 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10965 8144 6015 6103 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10964 7952 8171 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10963 8173 8172 7952 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10962 8144 8169 8173 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10961 2901 2690 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10960 2901 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10959 8144 4306 2901 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10958 165 3384 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10957 165 359 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10956 8144 1150 165 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10955 2674 3603 2676 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10954 2675 2887 2674 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10953 2673 2888 2675 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10952 8144 3606 2673 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10951 2672 2676 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10950 2215 2217 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10949 8144 5168 2215 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10948 2214 2215 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10947 2637 2847 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10946 8144 3229 2637 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10945 2642 2637 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10944 8144 7043 7036 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10943 7036 7034 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10942 8144 7038 7036 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10941 7033 7036 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10940 6307 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10939 6307 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10938 8144 6543 6307 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10937 8144 6076 6307 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10936 6340 6358 5996 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10935 5996 6359 6340 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10934 8144 7788 5996 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10933 5175 5445 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10932 8144 5178 5175 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10931 5642 5175 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10930 6137 7887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10929 6137 6138 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10928 8144 6161 6137 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10927 1986 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10926 1986 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10925 8144 4293 1986 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10924 4803 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10923 8144 7130 4803 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10922 344 166 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10921 344 365 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10920 8144 553 344 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10919 352 4251 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10918 352 359 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10917 8144 1150 352 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10916 2376 3780 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10915 8144 4255 2376 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10914 2375 2376 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10913 8144 3735 2603 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10912 2603 3730 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10911 8144 3744 2603 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10910 2601 2603 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10909 7062 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10908 7062 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10907 8144 6609 7062 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10906 8144 8097 7062 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10905 1372 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10904 1372 4067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10903 8144 5447 1372 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10902 8144 4228 1128 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10901 1128 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10900 1128 5147 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10899 8144 1372 1128 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10898 1788 1128 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10897 621 7548 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10896 765 764 621 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10895 620 1798 765 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10894 8144 1800 620 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10893 763 765 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10892 7251 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10891 7330 7798 7251 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10890 8144 7349 7330 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10889 5152 5151 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10888 8144 5154 5152 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10887 5150 5152 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10886 4695 5133 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10885 8144 4934 4695 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10884 4693 4695 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10883 2768 2890 2891 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10882 2766 7779 2768 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10881 2767 2889 2766 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10880 8144 7778 2767 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10879 3771 2891 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10878 1874 1905 2040 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10877 1875 2043 1874 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10876 8144 1904 1875 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10875 2041 2040 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10874 8144 6909 6419 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10873 6419 6636 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10872 8144 6921 6419 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10871 6418 6419 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10870 624 2968 777 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10869 625 5940 624 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10868 623 2262 625 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10867 8144 2964 623 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10866 778 777 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10865 2037 2036 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10864 8144 2035 2037 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10863 2485 2037 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10862 8144 2591 2593 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10861 2794 2589 2592 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10860 2592 2591 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10859 2592 2593 2794 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10858 8144 2590 2592 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10857 2590 2589 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10856 3510 5077 3509 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10855 8144 3507 3509 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10854 3509 7318 3510 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10853 3508 3510 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10852 8144 7398 6162 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10851 6162 7881 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10850 8144 8184 6162 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10849 6161 6162 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10848 6919 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10847 8144 7130 6919 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10846 7151 6919 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10845 1371 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10844 1370 4518 1371 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10843 1369 1372 1370 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10842 8144 2698 1369 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10841 1576 1370 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10840 5894 6273 5824 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10839 8144 5823 5824 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10838 5824 6480 5894 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10837 6051 5894 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10836 8144 5648 1830 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10835 1830 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10834 1830 5447 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10833 8144 7051 1830 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10832 1905 1830 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10831 8144 4051 4052 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10830 4052 4572 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10829 8144 5483 4052 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10828 4997 4052 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10827 986 1070 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10826 984 1072 1064 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10825 8144 1063 984 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10824 1072 1073 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10823 8144 1951 1073 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10822 8144 1069 1070 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10821 1067 1072 986 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10820 985 1073 1067 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10819 8144 1066 985 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10818 1066 1067 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10817 1064 1073 1066 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10816 8144 1064 1063 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10815 1063 1064 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10814 5851 5934 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10813 5849 5931 5930 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10812 8144 5938 5849 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10811 5931 5936 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10810 8144 7821 5936 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10809 8144 5935 5934 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10808 5933 5931 5851 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10807 5850 5936 5933 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10806 8144 5932 5850 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10805 5932 5933 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10804 5930 5936 5932 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10803 8144 5930 5938 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10802 5938 5930 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10801 7415 7750 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10800 7725 7747 7415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10799 8144 7793 7725 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10798 4728 4744 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10797 8144 4735 4728 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10796 3690 5453 4047 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10795 3689 8159 3690 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10794 8144 4734 3689 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10793 4030 5670 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10792 4556 4543 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10791 6304 5906 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10790 7750 7752 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10789 7766 7247 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10788 8046 7513 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10787 4213 5147 4088 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10786 8144 7802 4088 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10785 4088 5148 4213 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10784 4212 4213 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10783 910 912 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10782 906 914 907 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10781 8144 1317 906 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10780 914 913 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10779 8144 1772 913 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10778 8144 1074 912 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10777 911 914 910 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10776 908 913 911 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10775 8144 909 908 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10774 909 911 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10773 907 913 909 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10772 8144 907 1317 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10771 1317 907 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10770 8144 4995 4250 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10769 7871 4250 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10768 8144 4250 7871 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10767 8144 4250 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10766 8144 4250 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10765 8144 4995 4996 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10764 6383 4996 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10763 8144 4996 6383 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10762 8144 4996 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10761 8144 4996 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10760 8144 4552 4553 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10759 4995 4553 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10758 8144 4553 4995 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10757 8144 4553 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10756 8144 4553 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10755 8144 5616 5532 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10754 5532 6867 5617 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10753 5910 5617 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10752 7527 7788 7423 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10751 7423 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10750 8144 8021 7527 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10749 7525 7527 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10748 2752 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10747 4647 5907 2752 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10746 8144 6792 4647 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10745 1570 2492 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10744 8144 1799 1570 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10743 4009 6273 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10742 4413 6267 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10741 3716 6484 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10740 3602 5180 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10739 4933 5603 4931 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10738 4932 5906 4933 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10737 4933 6285 4932 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10736 4931 6286 4933 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10735 4931 6076 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10734 8144 6284 4931 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10733 1312 1738 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10732 4186 1739 1312 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10731 8144 3148 4186 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10730 3286 3100 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10729 8144 3095 3286 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10728 1297 1295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10727 1297 2168 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10726 8144 1296 1297 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10725 5076 5236 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10724 5074 5235 5229 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10723 8144 5227 5074 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10722 5235 5237 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10721 8144 5864 5237 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10720 8144 5232 5236 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10719 5234 5235 5076 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10718 5075 5237 5234 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10717 8144 5230 5075 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10716 5230 5234 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10715 5229 5237 5230 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10714 8144 5229 5227 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10713 5227 5229 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10712 6417 6917 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10711 8144 7140 6417 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10710 8169 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10709 8144 8159 8169 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10708 6402 6629 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10707 6401 6400 6402 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10706 8144 6399 6401 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10705 7550 2469 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10704 8144 4572 7550 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10703 1742 5830 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10702 8144 1741 1742 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10701 2176 4003 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10700 8144 2177 2176 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10699 2638 2176 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10698 2365 2166 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10697 8144 3229 2365 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10696 6434 6515 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10695 6432 6514 6508 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10694 8144 6506 6432 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10693 6514 6516 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10692 8144 8063 6516 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10691 8144 6513 6515 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10690 6510 6514 6434 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10689 6433 6516 6510 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10688 8144 6509 6433 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10687 6509 6510 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10686 6508 6516 6509 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10685 8144 6508 6506 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10684 6506 6508 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10683 7542 8097 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10682 7542 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10681 8144 7352 7542 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10680 5577 5576 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10679 8144 5574 5577 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10678 5897 5577 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10677 8144 7314 2926 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10676 8144 1807 1379 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10675 2926 1379 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10674 536 1115 538 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10673 538 1114 537 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10672 537 535 538 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10671 536 725 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10670 8144 1110 536 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10669 538 739 536 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10668 1965 537 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10667 5833 6300 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10666 8144 5905 5833 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10665 3114 3759 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10664 8144 4166 3114 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10663 5631 5628 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10662 8144 5629 5631 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10661 7747 5631 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10660 5637 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10659 5637 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10658 8144 5654 5637 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10657 8144 6375 5637 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10656 7106 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10655 7106 6909 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10654 8144 7880 7106 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10653 8144 7130 7106 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10652 6647 7398 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10651 8144 7891 6647 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10650 5840 6090 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10649 5917 6089 5840 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10648 8144 6567 5917 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10647 6466 4191 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10646 8144 4186 6466 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10645 1709 2132 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10644 1710 3737 1709 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10643 8144 2599 1710 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10642 2803 3586 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10641 2803 3293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10640 8144 3566 2803 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10639 8144 3581 2803 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10638 2856 3129 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_10637 2858 3135 2743 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10636 2743 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10635 8144 2854 2745 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10634 2745 2853 2744 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10633 2744 2856 2858 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10632 2858 3129 2746 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10631 2746 3145 2745 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10630 8144 3556 2854 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_10629 2860 2858 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10628 2650 3129 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_10627 2656 2648 2649 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10626 2649 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10625 8144 2651 2654 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10624 2654 2652 2653 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10623 2653 2650 2656 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10622 2656 3129 2655 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10621 2655 3143 2654 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10620 8144 3556 2651 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_10619 2873 2656 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10618 8144 6309 6310 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10617 6310 6307 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10616 8144 6308 6310 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10615 6536 6310 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10614 4596 6363 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10613 4719 4717 4596 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10612 4595 7343 4719 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10611 8144 4720 4595 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10610 5437 4719 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10609 8144 7091 7884 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10608 7091 7867 6940 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10607 6939 7094 7091 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10606 8144 7867 7094 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10605 6940 7549 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10604 8144 7272 6939 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10603 7884 7091 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10602 8144 5618 5431 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10601 5431 5620 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10600 5616 5428 5431 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10599 5430 5429 5616 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10598 5431 5432 5430 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10597 1427 5624 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10596 1538 4293 1427 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10595 8144 1992 1538 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10594 5970 5971 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10593 8144 8179 5970 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10592 6178 5970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10591 4253 7871 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10590 8144 4251 4253 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10589 4756 4253 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10588 5503 6172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10587 5503 6909 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10586 8144 7633 5503 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10585 8144 7130 5503 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10584 7701 7758 7757 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10583 7702 7787 7701 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10582 7700 8048 7702 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10581 8144 8045 7700 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10580 8004 7757 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10579 2700 4548 2701 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_10578 2699 2698 2700 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_10577 8144 5434 2699 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_10576 2701 2702 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_10575 5815 5881 7073 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10574 8144 7314 5881 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10573 5814 5888 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10572 7073 7314 5814 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10571 8144 5880 5815 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10570 3583 7343 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10569 3583 4228 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10568 8144 4517 3583 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10567 8144 4518 3583 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10566 8144 5648 3322 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10565 3322 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10564 3322 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10563 8144 6267 3322 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10562 3320 3322 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10561 4417 4914 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10560 4416 4502 4417 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10559 8144 4503 4416 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10558 6175 6909 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10557 8144 6172 6175 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10556 6407 6175 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10555 4899 5566 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10554 8144 5089 4899 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10553 4898 4899 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10552 157 163 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10551 156 159 157 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10550 155 342 156 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10549 8144 343 155 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10548 1115 156 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10547 8144 4538 4224 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10546 8144 4720 4223 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10545 4224 4223 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10544 5506 5718 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10543 8144 7352 5506 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10542 5505 5506 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10541 3157 3156 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10540 8144 3244 3157 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10539 3165 3157 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10538 998 1120 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10537 1122 1535 998 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10536 997 1541 1122 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10535 8144 1119 997 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10534 1785 1122 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10533 6483 6484 6424 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10532 8144 6481 6424 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10531 6424 6480 6483 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10530 6478 6483 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10529 6265 6267 6264 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10528 6264 6480 6265 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10527 8144 6266 6264 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10526 8144 7884 6660 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10525 6660 7892 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10524 6660 6893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10523 8144 7891 6660 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10522 6658 6660 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10521 8144 5453 5087 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10520 5384 5938 5046 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10519 5046 5453 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10518 5046 5087 5384 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10517 8144 5085 5046 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10516 5085 5938 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10515 8144 5863 4044 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10514 4044 8064 4045 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10513 8144 6797 2721 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10512 2721 6802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10511 2721 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10510 8144 3857 2721 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10509 2951 2721 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10508 3127 3763 3126 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10507 3126 4424 3127 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10506 8144 4510 3126 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10505 522 524 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10504 518 525 519 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10503 8144 517 518 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10502 525 526 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10501 8144 1772 526 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10500 8144 528 524 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10499 523 525 522 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10498 520 526 523 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10497 8144 521 520 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10496 521 523 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10495 519 526 521 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10494 8144 519 517 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10493 517 519 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10492 6368 6371 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10491 6365 6372 6366 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10490 8144 6602 6365 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10489 6372 6373 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10488 8144 7821 6373 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10487 8144 6600 6371 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10486 6369 6372 6368 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10485 6370 6373 6369 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10484 8144 6367 6370 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10483 6367 6369 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10482 6366 6373 6367 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10481 8144 6366 6602 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10480 6602 6366 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10479 5822 5891 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10478 5820 5892 5887 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10477 8144 5888 5820 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10476 5892 5893 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10475 8144 8063 5893 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10474 8144 7528 5891 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10473 5890 5892 5822 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10472 5821 5893 5890 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10471 8144 5889 5821 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10470 5889 5890 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10469 5887 5893 5889 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10468 8144 5887 5888 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10467 5888 5887 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10466 7785 7789 8028 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10465 7784 7782 7785 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10464 8144 7783 7784 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10463 8144 4472 4069 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10462 4072 4070 4074 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10461 4073 4315 4072 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10460 4069 4071 4073 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10459 78 79 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10458 74 80 73 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10457 8144 498 74 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10456 80 81 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10455 8144 1951 81 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10454 8144 261 79 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10453 76 80 78 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10452 77 81 76 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10451 8144 75 77 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10450 75 76 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10449 73 81 75 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10448 8144 73 498 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10447 498 73 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10446 6819 7257 7460 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10445 6818 6820 6819 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10444 8144 6816 6818 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10443 1303 1739 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10442 1473 1738 1303 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10441 8144 8045 1473 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10440 8144 4078 3655 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10439 3657 3667 3659 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10438 3658 3656 3657 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10437 3655 3851 3658 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10436 3687 3801 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10435 3802 4033 3687 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10434 8144 3804 3802 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10433 5008 5010 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10432 5004 5011 5005 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10431 8144 5003 5004 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10430 5011 5012 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10429 8144 5864 5012 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10428 8144 5226 5010 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10427 5009 5011 5008 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10426 5007 5012 5009 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10425 8144 5006 5007 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10424 5006 5009 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10423 5005 5012 5006 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10422 8144 5005 5003 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10421 5003 5005 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10420 1705 1707 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10419 1700 1706 1701 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10418 8144 5453 1700 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10417 1706 1708 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10416 8144 3708 1708 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10415 8144 2319 1707 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10414 1704 1706 1705 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10413 1703 1708 1704 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10412 8144 1702 1703 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10411 1702 1704 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10410 1701 1708 1702 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10409 8144 1701 5453 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10408 5453 1701 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10407 7310 7309 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10406 8144 7314 7310 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10405 8038 7772 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10404 8144 7773 8038 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10403 6188 5875 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10402 8144 6672 6188 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10401 7458 7321 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10400 8144 7322 7458 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10399 3553 3582 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10398 3553 3356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10397 8144 3581 3553 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10396 1455 3542 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10395 1455 3744 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10394 8144 2796 1455 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10393 1740 1739 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10392 2159 1738 1740 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10391 8144 1962 2159 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10390 5519 5614 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10389 5517 5613 5608 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10388 8144 5606 5517 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10387 5613 5615 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10386 8144 8063 5615 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10385 8144 5846 5614 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10384 5612 5613 5519 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10383 5518 5615 5612 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10382 8144 5609 5518 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10381 5609 5612 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10380 5608 5615 5609 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10379 8144 5608 5606 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10378 5606 5608 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10377 5161 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10376 5161 4224 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10375 8144 4310 5161 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10374 8144 6796 5161 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10373 6166 6636 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10372 6166 7121 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10371 8144 6652 6166 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10370 5908 5654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10369 5908 6609 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10368 8144 4302 5908 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10367 3851 3850 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10366 8144 4287 3851 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10365 2223 2688 2222 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10364 2222 2894 2221 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10363 2221 6796 2223 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10362 2223 2896 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10361 8144 4067 2223 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10360 2220 2221 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10359 2346 3348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10358 2346 3735 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10357 8144 3730 2346 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10356 2660 2661 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10355 2668 2659 2660 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10354 8144 2883 2668 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10353 4889 4892 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10352 4886 4893 4887 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10351 8144 6349 4886 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10350 4893 4894 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10349 8144 8063 4894 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10348 8144 5090 4892 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10347 4890 4893 4889 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10346 4891 4894 4890 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10345 8144 4888 4891 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10344 4888 4890 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10343 4887 4894 4888 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10342 8144 4887 6349 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10341 6349 4887 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10340 7522 7520 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10339 8144 7523 7522 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10338 7748 7522 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10337 4998 4999 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10336 4998 4997 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10335 8144 5000 4998 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10334 5712 5728 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10333 5712 6404 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10332 8144 5870 5712 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10331 6404 7887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10330 6404 6642 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10329 8144 6663 6404 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10328 3627 3625 3626 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10327 3626 6598 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10326 8144 3628 3627 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10325 3624 3627 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10324 8144 3788 3784 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10323 3784 3794 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10322 8144 4203 3784 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10321 3783 3784 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10320 2604 3293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10319 8144 3566 2604 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10318 2602 2604 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10317 3735 7585 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10316 3735 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10315 8144 4172 3735 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10314 8144 656 654 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10313 656 6867 585 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10312 584 658 656 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10311 8144 6867 658 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10310 585 3276 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10309 8144 6520 584 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10308 654 656 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10307 8144 4642 4641 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10306 4642 6867 4585 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10305 4584 4645 4642 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10304 8144 6867 4645 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10303 4585 4644 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10302 8144 6292 4584 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10301 4641 4642 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10300 8144 3960 3955 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10299 3960 6867 3959 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10298 3957 3961 3960 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10297 8144 6867 3961 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10296 3959 3958 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10295 8144 3956 3957 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10294 3955 3960 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10293 8144 3618 3383 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10292 3383 3378 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10291 8144 3379 3383 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10290 5426 3383 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10289 5498 5868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10288 5498 5971 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10287 8144 7633 5498 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10286 1801 1800 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10285 3170 1798 1801 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10284 8144 3150 3170 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10283 349 4558 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10282 349 359 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10281 8144 1150 349 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10280 8144 3966 3962 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10279 3966 6867 3965 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10278 3963 3967 3966 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10277 8144 6867 3967 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10276 3965 3964 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10275 8144 6792 3963 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10274 3962 3966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10273 6554 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10272 6554 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10271 8144 7026 6554 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10270 8144 6080 6554 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10269 7436 7563 7591 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10268 8144 7957 7563 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10267 7435 7835 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10266 7591 7957 7435 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10265 8144 7970 7436 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10264 5373 5880 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10263 8144 7500 5373 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10262 7708 8009 7771 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10261 7707 7787 7708 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10260 7706 8048 7707 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10259 8144 8045 7706 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10258 7773 7771 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10257 5047 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10256 5089 5907 5047 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10255 8144 6349 5089 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10254 3696 4734 3837 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10253 3695 5453 3696 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10252 8144 8159 3695 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10251 3839 3837 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10250 6270 6485 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10249 8144 7500 6270 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10248 4513 4932 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10247 8144 4953 4513 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10246 4427 4513 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10245 8144 7881 7394 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10244 7394 7408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10243 8144 7883 7394 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10242 7872 7394 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10241 3713 4130 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10240 8144 3714 3713 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10239 3711 3713 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10238 3678 4413 3724 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10237 3676 7787 3678 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10236 3677 8048 3676 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10235 8144 8045 3677 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10234 3723 3724 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10233 6952 7065 7612 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10232 8144 7957 7065 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10231 6953 7558 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10230 7612 7957 6953 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10229 8144 7803 6952 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10228 3778 5147 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10227 8144 5148 3778 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10226 3776 3778 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10225 162 365 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10224 8144 166 162 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10223 161 162 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10222 1844 4189 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10221 1954 2170 1844 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10220 8144 2375 1954 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10219 8144 7398 6645 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10218 6645 7892 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10217 8144 7869 6645 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10216 6642 6645 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10215 8144 4896 4897 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10214 4897 4902 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10213 8144 5606 4897 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10212 4895 4897 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10211 8144 2719 1828 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10210 1828 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10209 8144 3857 1828 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10208 1827 1828 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10207 8144 7881 6405 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10206 6405 6893 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10205 8144 7891 6405 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10204 6636 6405 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10203 102 101 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10202 97 103 96 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10201 8144 273 97 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10200 103 104 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10199 8144 1951 104 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10198 8144 272 101 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10197 100 103 102 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10196 98 104 100 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10195 8144 99 98 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10194 99 100 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10193 96 104 99 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10192 8144 96 273 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10191 273 96 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10190 8144 7247 7311 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10189 8144 7957 6762 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10188 7311 6762 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10187 8144 4068 3815 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10186 3815 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10185 8144 4574 3815 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10184 3812 3815 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10183 8144 6802 958 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10182 958 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10181 958 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10180 8144 6796 958 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10179 1167 958 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10178 5417 6506 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10177 4406 6489 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10176 4705 6775 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10175 1419 1956 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10174 2361 1957 1419 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10173 8144 1962 2361 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10172 2835 3112 2755 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10171 2755 3111 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10170 8144 3108 2835 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10169 2833 2835 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10168 5473 5475 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10167 5469 5477 5470 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10166 8144 5664 5469 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10165 5477 5476 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10164 8144 5864 5476 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10163 8144 5478 5475 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10162 5474 5477 5473 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10161 5472 5476 5474 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10160 8144 5471 5472 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10159 5471 5474 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10158 5470 5476 5471 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10157 8144 5470 5664 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10156 5664 5470 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10155 5896 5394 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10154 5896 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10153 8144 7352 5896 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10152 5111 5113 5052 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10151 5052 5118 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10150 8144 5110 5111 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10149 5109 5111 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_10148 3252 3623 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10147 8144 4048 3252 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10146 4999 5202 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10145 6594 6602 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10144 4260 5227 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10143 4032 4760 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10142 5429 5603 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10141 5413 5898 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10140 1404 1508 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10139 1402 1507 1501 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10138 8144 1499 1402 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10137 1507 1509 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10136 8144 1772 1509 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10135 8144 1506 1508 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10134 1504 1507 1404 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10133 1403 1509 1504 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10132 8144 1502 1403 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10131 1502 1504 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10130 1501 1509 1502 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10129 8144 1501 1499 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10128 1499 1501 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10127 4096 4268 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10126 4094 4267 4262 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10125 8144 4770 4094 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10124 4267 4269 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10123 8144 5864 4269 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10122 8144 4769 4268 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10121 4266 4267 4096 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10120 4095 4269 4266 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10119 8144 4263 4095 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10118 4263 4266 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10117 4262 4269 4263 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10116 8144 4262 4770 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10115 4770 4262 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10114 7914 8036 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10113 7912 8035 8030 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10112 8144 8040 7912 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10111 8035 8037 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10110 8144 8063 8037 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10109 8144 8039 8036 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10108 8034 8035 7914 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10107 7913 8037 8034 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10106 8144 8031 7913 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10105 8031 8034 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10104 8030 8037 8031 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10103 8144 8030 8040 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10102 8040 8030 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10101 6298 5419 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10100 6298 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10099 8144 7352 6298 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10098 1798 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10097 8144 5942 1798 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10096 6524 6292 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10095 8144 1616 1388 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10094 1391 1389 2035 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10093 1392 1390 1391 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10092 1388 1615 1392 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10091 2502 4427 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10090 8144 2172 2502 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10089 7243 7318 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10088 7309 7503 7243 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10087 8144 7316 7309 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10086 956 3608 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10085 8144 957 956 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10084 951 946 952 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10083 949 947 951 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10082 950 1139 949 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10081 8144 948 950 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_10080 1119 952 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10079 5241 5502 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10078 8144 5724 5241 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10077 6128 5944 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10076 8144 6137 6128 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10075 5944 5937 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10074 8144 6127 5944 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10073 7882 7881 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10072 8144 7891 7882 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10071 7453 7643 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10070 7646 8186 7453 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10069 8144 7869 7646 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10068 8144 2968 626 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10067 627 5940 2719 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10066 628 2262 627 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10065 626 2964 628 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10064 3580 3780 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10063 8144 5197 3580 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10062 3579 3580 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10061 5513 5583 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10060 5511 5585 5579 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10059 8144 5898 5511 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10058 5585 5586 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10057 8144 8063 5586 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_10056 8144 5589 5583 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10055 5582 5585 5513 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10054 5512 5586 5582 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10053 8144 5580 5512 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10052 5580 5582 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10051 5579 5586 5580 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_10050 8144 5579 5898 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10049 5898 5579 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10048 6309 6080 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10047 6309 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10046 8144 7352 6309 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10045 5468 5682 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10044 8144 5665 5468 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_10043 5467 5468 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10042 8144 7371 7271 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10041 7371 8140 7274 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10040 7273 7275 7371 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10039 8144 8140 7275 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10038 7274 7549 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10037 8144 7272 7273 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10036 7271 7371 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10035 8144 7375 7575 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10034 7375 8140 7277 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10033 7276 7278 7375 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10032 8144 8140 7278 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10031 7277 7528 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10030 8144 7572 7276 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10029 7575 7375 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10028 8144 7579 7851 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10027 7579 8140 7440 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10026 7439 7580 7579 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10025 8144 8140 7580 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10024 7440 7585 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10023 8144 7845 7439 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10022 7851 7579 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10021 8144 7386 7384 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10020 7386 8140 7288 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10019 7287 7289 7386 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10018 8144 8140 7289 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10017 7288 7349 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10016 8144 7379 7287 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10015 7384 7386 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10014 8144 7606 7603 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10013 7606 8140 7448 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10012 7447 7608 7606 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10011 8144 8140 7608 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10010 7448 7777 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10009 8144 7604 7447 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10008 7603 7606 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10007 8144 6852 6907 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10006 6852 7867 6851 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10005 6849 6853 6852 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10004 8144 7867 6853 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10003 6851 6850 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10002 8144 7076 6849 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_10001 6907 6852 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_10000 3542 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09999 3542 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09998 8144 4574 3542 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09997 8144 6484 3542 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09996 8144 8142 8153 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09995 8142 8140 7945 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09994 7944 8143 8142 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09993 8144 8140 8143 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09992 7945 8139 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09991 8144 8147 7944 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09990 8153 8142 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09989 8144 7861 8130 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09988 7861 8140 7720 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09987 7719 7862 7861 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09986 8144 8140 7862 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09985 7720 7863 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09984 8144 8125 7719 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09983 8130 7861 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09982 5491 6629 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09981 5490 5866 5491 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09980 8144 5489 5490 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09979 4317 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09978 4317 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09977 8144 4575 4317 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09976 8144 5483 4317 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09975 7249 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09974 7322 7798 7249 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09973 8144 7528 7322 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09972 1936 1943 1415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09971 1415 2154 1936 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09970 8144 2616 1415 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09969 3566 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09968 3566 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09967 8144 4167 3566 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09966 8144 6267 3566 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09965 8144 5574 4710 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09964 4710 5434 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09963 8144 6363 4710 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09962 4707 4710 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09961 8144 2203 2204 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09960 2204 7343 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09959 2204 5148 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09958 8144 4548 2204 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09957 4172 2204 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09956 8144 5673 5671 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09955 5673 6383 5522 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09954 5523 5675 5673 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09953 8144 6383 5675 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09952 5522 5858 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09951 8144 5670 5523 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09950 5671 5673 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09949 8144 7600 7643 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09948 7600 7867 7446 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09947 7445 7601 7600 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09946 8144 7867 7601 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09945 7446 7863 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09944 8144 8125 7445 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09943 7643 7600 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09942 8144 1788 1789 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09941 1789 2214 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09940 1789 1985 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09939 8144 2207 1789 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09938 4173 1789 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09937 6283 6784 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09936 6502 6785 6283 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09935 8144 7500 6502 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09934 6962 7304 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09933 7400 7151 6962 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09932 8144 7149 7400 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09931 6154 6158 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09930 6154 6157 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09929 8144 6156 6154 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09928 8144 6166 6154 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09927 8144 5120 4696 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09926 4698 7059 4592 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09925 4592 5120 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09924 4592 4696 4698 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09923 8144 4697 4592 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09922 4697 7059 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09921 6766 7559 6764 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09920 6764 7548 6765 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09919 6765 7550 6766 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09918 6766 6972 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09917 8144 6985 6766 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09916 6763 6765 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09915 4409 4406 4490 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09914 4407 7787 4409 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09913 4408 8048 4407 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09912 8144 8045 4408 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09911 4405 4490 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09910 1316 1956 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09909 1315 1957 1316 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09908 8144 8045 1315 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09907 2466 1816 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09906 2466 1817 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09905 8144 1818 2466 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09904 8144 1819 2466 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09903 1314 1957 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09902 1313 1956 1314 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09901 8144 3148 1313 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09900 8144 865 860 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09899 3276 2595 859 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09898 859 865 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09897 859 860 3276 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09896 8144 858 859 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09895 858 2595 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09894 7419 8046 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09893 7518 7747 7419 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09892 8144 7517 7518 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09891 7549 6850 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09890 4066 5032 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09889 8144 4790 4066 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09888 4071 4066 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09887 1329 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09886 8144 1335 1329 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09885 1327 1329 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09884 4105 7056 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09883 4183 5406 4105 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09882 8144 6812 4183 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09881 6782 6781 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09880 6780 6778 6782 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09879 8144 6779 6780 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09878 8144 7881 5969 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09877 5969 8187 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09876 8144 7883 5969 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09875 5971 5969 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09874 769 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09873 8144 5483 769 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09872 1140 769 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09871 8144 2234 2237 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09870 2237 2235 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09869 8144 2236 2237 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09868 2246 2237 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09867 5847 6375 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09866 6325 5922 5847 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09865 8144 5923 6325 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09864 8144 4803 4806 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09863 4806 4802 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09862 8144 5044 4806 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09861 4801 4806 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09860 1756 1965 1757 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09859 1757 1964 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09858 8144 1962 1756 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09857 2174 1756 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09856 1848 2178 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09855 3128 2179 1848 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09854 8144 1962 3128 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09853 136 138 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09852 132 139 133 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09851 8144 530 132 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09850 139 140 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09849 8144 1772 140 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09848 8144 141 138 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09847 137 139 136 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09846 135 140 137 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09845 8144 134 135 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09844 134 137 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09843 133 140 134 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09842 8144 133 530 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09841 530 133 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09840 8144 558 358 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09839 358 559 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09838 358 1362 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09837 8144 6363 358 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09836 359 358 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09835 600 1115 601 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09834 601 1114 708 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09833 708 709 601 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09832 600 703 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09831 8144 1110 600 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09830 601 900 600 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09829 1957 708 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09828 1006 1116 1005 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09827 1348 1113 1006 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09826 1006 1114 1348 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09825 1005 1115 1006 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09824 1005 1111 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09823 8144 1110 1005 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09822 1930 2595 1838 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09821 1838 2138 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09820 8144 1929 1930 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09819 1928 1930 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09818 195 197 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09817 191 198 192 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09816 8144 190 191 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09815 198 199 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09814 8144 3834 199 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09813 8144 1699 197 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09812 196 198 195 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09811 194 199 196 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09810 8144 193 194 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09809 193 196 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09808 192 199 193 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09807 8144 192 190 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09806 190 192 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09805 6928 6981 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09804 6926 6982 6976 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09803 8144 6974 6926 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09802 6982 6983 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09801 8144 8063 6983 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09800 8144 7585 6981 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09799 6979 6982 6928 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09798 6927 6983 6979 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09797 8144 6977 6927 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09796 6977 6979 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09795 6976 6983 6977 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09794 8144 6976 6974 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09793 6974 6976 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09792 7921 8053 8067 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09791 7920 8054 7921 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09790 8144 8052 7920 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09789 6950 7056 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09788 7359 7058 6950 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09787 8144 7342 7359 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09786 8144 4295 1385 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09785 1385 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09784 1385 4167 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09783 8144 5624 1385 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09782 1384 1385 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09781 3612 4032 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09780 3611 3610 3612 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09779 8144 3613 3611 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09778 616 753 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09777 614 752 747 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09776 8144 1116 614 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09775 752 754 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09774 8144 3834 754 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09773 8144 751 753 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09772 748 752 616 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09771 615 754 748 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09770 8144 749 615 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09769 749 748 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09768 747 754 749 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09767 8144 747 1116 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09766 1116 747 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09765 6461 6626 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09764 6459 6625 6620 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09763 8144 6618 6459 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09762 6625 6628 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09761 8144 8166 6628 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09760 8144 6630 6626 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09759 6624 6625 6461 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09758 6460 6628 6624 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09757 8144 6622 6460 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09756 6622 6624 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09755 6620 6628 6622 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09754 8144 6620 6618 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09753 6618 6620 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09752 4091 4247 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09751 4089 4248 4241 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09750 8144 4955 4089 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09749 4248 4249 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09748 8144 5864 4249 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09747 8144 4244 4247 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09746 4245 4248 4091 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09745 4090 4249 4245 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09744 8144 4242 4090 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09743 4242 4245 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09742 4241 4249 4242 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09741 8144 4241 4955 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09740 4955 4241 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09739 215 3956 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09738 8144 3956 241 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09737 238 2127 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09736 8144 238 215 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09735 215 241 240 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09734 240 2127 215 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09733 1446 240 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09732 8144 240 1446 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09731 8144 6921 6414 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09730 6414 7148 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09729 6412 7151 6414 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09728 6413 6655 6412 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09727 6414 6658 6413 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09726 8066 8028 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09725 8144 8025 8066 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09724 7556 7788 7434 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09723 7434 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09722 8144 8071 7556 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09721 8053 7556 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09720 2316 5633 2272 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09719 2272 2789 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09718 8144 5372 2316 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09717 2315 2316 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09716 4578 5245 4469 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09715 4469 4583 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09714 8144 4577 4578 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09713 4468 4578 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09712 3587 4203 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09711 3587 3788 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09710 8144 3794 3587 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09709 3737 3582 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09708 3737 3356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09707 8144 3579 3737 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09706 8144 3744 2137 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09705 2137 2135 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09704 2133 2599 2137 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09703 2134 2132 2133 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09702 2137 3737 2134 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09701 854 855 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09700 849 856 850 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09699 8144 2127 849 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09698 856 857 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09697 8144 3708 857 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09696 8144 2126 855 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09695 853 856 854 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09694 852 857 853 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09693 8144 851 852 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09692 851 853 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09691 850 857 851 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09690 8144 850 2127 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09689 2127 850 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09688 7147 8184 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09687 7147 7403 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09686 8144 7884 7147 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09685 8089 7460 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09684 8144 7801 8089 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09683 4078 4474 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09682 8144 4477 4078 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09681 2242 2027 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09680 2242 2448 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09679 8144 2251 2242 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09678 4964 4965 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09677 4959 4967 4958 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09676 8144 6341 4959 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09675 4967 4966 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09674 8144 7821 4966 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09673 8144 4963 4965 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09672 4961 4967 4964 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09671 4962 4966 4961 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09670 8144 4960 4962 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09669 4960 4961 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09668 4958 4966 4960 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09667 8144 4958 6341 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09666 6341 4958 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09665 4908 4910 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09664 4904 4911 4905 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09663 8144 6801 4904 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09662 4911 4912 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09661 8144 8063 4912 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09660 8144 4913 4910 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09659 4909 4911 4908 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09658 4907 4912 4909 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09657 8144 4906 4907 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09656 4906 4909 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09655 4905 4912 4906 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09654 8144 4905 6801 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09653 6801 4905 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09652 5527 6793 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09651 6266 6294 5527 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09650 8144 5553 6266 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09649 5165 5161 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09648 8144 5160 5165 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09647 5162 5165 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09646 1786 1790 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09645 8094 1785 1786 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09644 8144 7314 8094 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09643 6470 7730 6423 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09642 6423 7738 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09641 8144 8064 6470 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09640 6469 6470 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09639 3604 3611 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09638 8144 6341 3604 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09637 3603 3604 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09636 1300 1476 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09635 1466 1477 1300 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09634 8144 1962 1466 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09633 5126 5164 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09632 8144 7012 5126 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09631 5124 5126 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09630 8144 4917 4913 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09629 4917 6867 4915 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09628 4916 4918 4917 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09627 8144 6867 4918 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09626 4915 4914 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09625 8144 6801 4916 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09624 4913 4917 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09623 8144 5094 5090 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09622 5094 6867 5049 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09621 5048 5095 5094 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09620 8144 6867 5095 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09619 5049 5092 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09618 8144 6349 5048 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09617 5090 5094 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09616 6262 6786 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09615 6262 6051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09614 8144 6500 6262 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09613 8144 6503 6262 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09612 5870 5968 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09611 5870 6909 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09610 8144 6921 5870 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09609 760 1353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09608 760 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09607 8144 5483 760 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09606 8144 2202 1694 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09605 1694 2199 1775 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09604 1776 1775 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09603 8144 4509 4681 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09602 4509 6867 4421 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09601 4422 4423 4509 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09600 8144 6867 4423 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09599 4421 4502 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09598 8144 6549 4422 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09597 4681 4509 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09596 8144 7542 7546 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09595 7546 7541 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09594 8144 7543 7546 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09593 7794 7546 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09592 8144 6478 4118 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09591 4118 6472 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09590 8144 6473 4118 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09589 5078 4118 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09588 8144 6786 6281 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09587 6281 6500 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09586 6281 6784 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09585 8144 6785 6281 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09584 6778 6281 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09583 8144 6618 6335 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09582 8144 6549 6018 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09581 6335 6018 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09580 7395 7300 7298 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09579 8144 7871 7298 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09578 7298 7875 7395 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09577 7297 7395 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09576 6671 6670 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09575 8144 7405 6671 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09574 6668 6671 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09573 5728 6921 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09572 5728 6176 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09571 8144 5875 5728 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09570 8144 1807 1011 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09569 1011 8064 1160 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09568 2698 1160 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09567 8144 8159 2777 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09566 2777 5453 2923 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09565 2922 2923 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09564 8144 5940 2261 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09563 2260 2261 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09562 8144 2262 2260 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09561 2490 2260 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09560 8144 2260 2490 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09559 6532 6804 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09558 8144 7500 6532 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09557 1987 7559 1854 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09556 1854 7548 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09555 8144 1986 1987 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09554 2205 1987 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09553 1413 3737 1412 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09552 1412 2132 1453 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09551 1453 2599 1413 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09550 1413 2135 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09549 8144 3744 1413 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09548 1451 1453 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09547 8144 4167 3727 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09546 3727 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09545 3727 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09544 8144 6273 3727 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09543 3725 3727 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09542 6439 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09541 6540 7798 6439 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09540 8144 8122 6540 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09539 5966 6409 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09538 8144 5967 5966 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09537 5869 5966 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09536 7919 8046 8049 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09535 7917 8047 7919 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09534 7918 8048 7917 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09533 8144 8045 7918 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09532 8068 8049 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09531 4470 4790 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09530 4470 6421 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09529 8144 6672 4470 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09528 8144 5740 4470 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09527 6972 6987 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09526 8144 7957 6972 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09525 8144 6359 1994 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09524 1994 1887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09523 1994 2924 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09522 8144 1891 1994 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09521 2207 1994 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09520 6795 6793 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09519 7459 7058 6795 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09518 8144 6794 7459 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09517 5914 5912 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09516 8144 5913 5914 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09515 5837 5914 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09514 7804 7803 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09513 8144 7957 7804 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09512 5973 7408 5877 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09511 5877 7893 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09510 8144 8184 5973 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09509 5876 5973 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09508 4799 5034 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09507 8144 4801 4799 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09506 4798 4799 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09505 3879 3877 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09504 8144 4318 3879 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09503 3876 3879 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09502 2208 7343 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09501 8144 2227 2208 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09500 2421 2208 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09499 4426 4511 4425 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09498 4425 4512 4426 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09497 8144 4510 4425 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09496 8144 7884 6911 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09495 6911 7403 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09494 6911 7408 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09493 8144 8184 6911 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09492 6917 6911 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09491 1305 5641 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09490 8144 1304 1305 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09489 1739 1305 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09488 2341 3725 2280 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09487 2280 2614 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09486 8144 3315 2341 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09485 2340 2341 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09484 7487 7486 7410 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09483 8144 7484 7410 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09482 7410 7490 7487 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09481 7485 7487 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09480 8144 6311 3401 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09479 3401 4573 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09478 8144 4293 3401 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09477 3844 3401 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09476 8144 3260 3418 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09475 3418 3659 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09474 3418 3858 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09473 8144 3261 3418 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09472 3419 3418 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09471 8144 3794 3149 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09470 3149 4203 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09469 8144 5908 3149 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09468 3148 3149 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09467 8144 7314 1450 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09466 1448 1450 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09465 8144 6267 1448 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09464 6084 1448 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09463 8144 1448 6084 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09462 6457 6870 6607 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09461 6456 7095 6457 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09460 8144 6618 6456 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09459 8144 6609 3617 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09458 3617 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09457 8144 5447 3617 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09456 3809 3617 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09455 8144 3416 3181 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09454 3181 3182 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09453 8144 3410 3181 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09452 3187 3181 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09451 8144 4293 2259 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09450 2259 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09449 2259 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09448 8144 5654 2259 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09447 2258 2259 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09446 8144 5265 5258 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09445 5258 5505 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09444 5258 5730 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09443 8144 5262 5258 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09442 5256 5258 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09441 8144 6185 5035 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09440 5035 5040 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09439 5035 5256 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09438 8144 5036 5035 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09437 5034 5035 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09436 597 693 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09435 595 692 684 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09434 8144 685 595 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09433 692 694 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09432 8144 1951 694 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09431 8144 691 693 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09430 686 692 597 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09429 596 694 686 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09428 8144 688 596 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09427 688 686 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09426 684 694 688 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09425 8144 684 685 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09424 685 684 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09423 4040 4041 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09422 4035 4042 4036 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09421 8144 4255 4035 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09420 4042 4043 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09419 8144 5864 4043 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09418 8144 4254 4041 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09417 4039 4042 4040 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09416 4038 4043 4039 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09415 8144 4037 4038 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09414 4037 4039 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09413 4036 4043 4037 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09412 8144 4036 4255 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09411 4255 4036 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09410 6793 6520 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09409 4896 5453 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09408 7020 6792 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09407 6821 6541 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09406 7029 6349 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09405 7056 6801 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09404 8144 2254 2253 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09403 2253 2252 3184 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09402 8144 4688 3684 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09401 3684 3997 3758 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09400 3757 3758 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09399 3119 3575 3120 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09398 3120 3121 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09397 8144 3118 3119 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09396 3310 3119 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09395 606 721 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09394 604 722 715 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09393 8144 1088 604 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09392 722 723 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09391 8144 1772 723 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09390 8144 915 721 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09389 716 722 606 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09388 605 723 716 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09387 8144 718 605 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09386 718 716 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09385 715 723 718 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09384 8144 715 1088 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09383 1088 715 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09382 5576 5571 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09381 5576 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09380 8144 7041 5576 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09379 4443 4538 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09378 4717 4530 4443 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09377 8144 5443 4717 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09376 5842 5908 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09375 8144 6363 5842 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09374 7531 7778 7424 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09373 7424 7779 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09372 8144 7528 7531 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09371 7529 7531 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09370 2241 2236 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09369 2241 2234 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09368 8144 2235 2241 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09367 8144 1169 1017 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09366 1015 1173 2247 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09365 1016 1167 1015 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09364 1017 1168 1016 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09363 3251 2912 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09362 8144 2913 3251 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09361 4901 5108 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09360 4902 5938 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09359 7059 6549 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09358 4939 6076 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09357 8144 2249 1869 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09356 1870 1898 2484 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09355 1868 2454 1870 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09354 1869 1897 1868 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09353 2594 2591 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09352 8144 2143 2594 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09351 7928 8082 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09350 7926 8083 8077 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09349 8144 8086 7926 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09348 8083 8084 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09347 8144 8166 8084 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09346 8144 8085 8082 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09345 8079 8083 7928 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09344 7927 8084 8079 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09343 8144 8078 7927 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09342 8078 8079 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09341 8077 8084 8078 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09340 8144 8077 8086 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09339 8086 8077 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09338 8144 1352 1354 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09337 1354 1353 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09336 1539 2210 1354 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09335 1351 5624 1539 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09334 1354 4293 1351 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09333 5935 6132 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09332 8144 5939 5935 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09331 4525 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09330 4525 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09329 8144 7354 4525 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09328 4540 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09327 4540 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09326 8144 6311 4540 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09325 1571 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09324 8144 4574 1571 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09323 2689 4293 2686 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09322 2686 4067 2685 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09321 2685 3370 2689 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09320 2689 2687 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09319 8144 2688 2689 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09318 7778 2685 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09317 1949 4685 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09316 8144 2361 1949 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09315 2352 1949 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09314 5516 5598 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09313 5514 5597 5592 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09312 8144 5603 5514 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09311 5597 5599 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09310 8144 8063 5599 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09309 8144 5835 5598 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09308 5594 5597 5516 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09307 5515 5599 5594 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09306 8144 5593 5515 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09305 5593 5594 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09304 5592 5599 5593 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09303 8144 5592 5603 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09302 5603 5592 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09301 6075 6554 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09300 8144 7343 6075 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09299 6308 6075 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09298 5561 5562 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09297 8144 7343 5561 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09296 5886 5561 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09295 8144 8121 8118 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09294 8121 8140 7940 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09293 7939 8124 8121 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09292 8144 8140 8124 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09291 7940 8122 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09290 8144 8119 7939 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09289 8118 8121 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09288 5939 5937 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09287 8144 5938 5939 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09286 2203 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09285 2203 1565 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09284 8144 6609 2203 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09283 2227 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09282 2227 1565 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09281 8144 6802 2227 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09280 1745 1744 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09279 5905 1743 1745 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09278 8144 3148 5905 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09277 2336 3735 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09276 8144 3730 2336 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09275 2334 2336 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09274 8144 5184 5181 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09273 5184 7871 5059 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09272 5060 5185 5184 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09271 8144 7871 5185 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09270 5059 5693 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09269 8144 5180 5060 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09268 5181 5184 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09267 4552 7353 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09266 4552 5654 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09265 8144 5483 4552 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09264 8144 7500 4552 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09263 8144 7345 6803 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09262 8144 7957 6805 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09261 6803 6805 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09260 8144 1807 962 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09259 961 962 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09258 8144 7314 961 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09257 963 961 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09256 8144 961 963 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09255 8144 7856 7888 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09254 7856 7867 7716 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09253 7715 7857 7856 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09252 8144 7867 7857 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09251 7716 8058 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09250 8144 7858 7715 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09249 7888 7856 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09248 8144 7859 8186 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09247 7859 7867 7718 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09246 7717 7860 7859 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09245 8144 7867 7860 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09244 7718 8122 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09243 8144 8119 7717 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09242 8186 7859 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09241 8144 7590 7619 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09240 7590 7867 7444 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09239 7443 7593 7590 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09238 8144 7867 7593 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09237 7444 7591 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09236 8144 7596 7443 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09235 7619 7590 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09234 8144 2006 1862 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09233 1862 2707 2010 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09232 2011 2010 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09231 8144 3819 1360 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09230 1360 1358 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09229 8144 1359 1360 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09228 1357 1360 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09227 2611 2614 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09226 2610 3725 2611 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09225 8144 3315 2610 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09224 8144 3744 3101 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09223 3101 3104 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09222 3100 3102 3101 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09221 3099 3737 3100 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09220 3101 3098 3099 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09219 2640 2648 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_09218 2646 2638 2639 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09217 2639 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09216 8144 2641 2644 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09215 2644 2642 2643 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09214 2643 2640 2646 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09213 2646 2648 2645 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09212 2645 3330 2644 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09211 8144 3556 2641 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_09210 3567 2646 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09209 8144 6974 6271 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09208 8144 7500 6272 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09207 6271 6272 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09206 8144 7614 7630 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09205 7614 7867 7450 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09204 7449 7615 7614 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09203 8144 7867 7615 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09202 7450 7612 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09201 8144 8137 7449 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09200 7630 7614 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09199 8144 7865 8187 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09198 7865 7867 7722 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09197 7721 7866 7865 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09196 8144 7867 7866 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09195 7722 8139 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09194 8144 8147 7721 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09193 8187 7865 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09192 8144 4574 3994 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09191 3994 7356 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09190 3994 6293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09189 8144 6775 3994 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09188 3993 3994 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09187 2621 2827 2281 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09186 2281 3307 2621 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09185 8144 2616 2281 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09184 2384 2648 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_09183 2387 2379 2292 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09182 2292 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09181 8144 2380 2295 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09180 2295 2382 2293 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09179 2293 2384 2387 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09178 2387 2648 2294 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09177 2294 3127 2295 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09176 8144 3556 2380 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_09175 2845 2387 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09174 3512 4885 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09173 3511 5078 3512 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09172 8144 3765 3511 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09171 8144 8176 7397 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09170 7397 7399 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09169 8144 7400 7397 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09168 7300 7397 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09167 8144 2202 1779 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09166 1777 1779 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09165 8144 1780 1777 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09164 1778 1777 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09163 8144 1777 1778 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09162 7704 7766 7764 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09161 7705 7787 7704 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09160 7703 8048 7705 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09159 8144 8045 7703 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09158 7765 7764 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09157 6289 6489 6287 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09156 6288 7513 6289 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09155 6289 6285 6288 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09154 6287 6286 6289 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09153 6287 6349 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09152 8144 6284 6287 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09151 7501 7742 7413 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09150 7413 7754 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09149 8144 7500 7501 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09148 7741 7501 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09147 2291 2840 2290 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09146 2290 2379 2373 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09145 2373 2371 2291 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09144 2291 4255 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09143 8144 3780 2291 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09142 2631 2373 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09141 8144 2794 2795 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09140 3964 3287 2753 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09139 2753 2794 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09138 2753 2795 3964 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09137 8144 2791 2753 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09136 2791 3287 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09135 8144 6506 6504 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09134 8144 7957 6282 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09133 6504 6282 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09132 2807 2806 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09131 8144 3723 2807 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09130 2805 2807 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09129 1349 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09128 8144 7026 1349 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09127 2210 1349 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09126 4742 4734 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09125 5178 5664 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09124 6867 7957 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09123 4739 5863 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09122 6586 6870 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09121 3843 3839 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09120 8144 4075 3843 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09119 3841 3843 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09118 8144 2132 862 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09117 862 1451 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09116 1292 1929 862 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09115 861 1287 1292 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09114 862 2595 861 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09113 6086 6087 5991 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09112 8144 6084 5991 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09111 5991 6083 6086 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_09110 6085 6086 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09109 6296 6821 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09108 6295 6294 6296 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09107 8144 6297 6295 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09106 2230 2926 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09105 2228 5148 2230 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09104 2229 4518 2228 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09103 8144 2698 2229 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09102 2236 2228 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09101 3183 3182 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09100 8144 3410 3183 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09099 3261 3183 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09098 4722 4720 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09097 4731 4538 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09096 6142 6141 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09095 6358 6618 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09094 6381 6143 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09093 8144 161 158 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09092 158 165 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09091 158 551 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09090 8144 349 158 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09089 1114 158 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09088 5982 6484 5981 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09087 6062 7979 5982 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09086 5982 6285 6062 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09085 5981 6286 5982 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09084 5981 6292 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09083 8144 6284 5981 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09082 7739 7802 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09081 7738 7747 7739 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09080 8144 7737 7738 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09079 8144 8064 2788 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09078 2787 2788 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09077 8144 5906 2787 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09076 3507 2787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09075 8144 2787 3507 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09074 1783 7559 1784 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09073 1784 7548 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09072 8144 1891 1783 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09071 1782 1783 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_09070 2684 2894 2681 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09069 2681 2898 2683 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09068 2683 4067 2684 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09067 2684 2682 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09066 8144 6796 2684 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09065 7779 2683 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09064 8144 6802 1595 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09063 1595 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09062 1595 6543 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09061 8144 5624 1595 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09060 1597 1595 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09059 8144 8159 3691 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09058 3691 5453 3826 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09057 8144 6543 4278 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09056 4278 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09055 4278 5942 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09054 8144 7051 4278 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09053 4280 4278 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09052 3750 1297 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09051 8144 1298 3750 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_09050 172 174 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09049 168 175 169 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09048 8144 4538 168 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09047 175 176 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09046 8144 3834 176 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09045 8144 177 174 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09044 173 175 172 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09043 171 176 173 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09042 8144 170 171 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09041 170 173 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09040 169 176 170 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09039 8144 169 4538 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09038 4538 169 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09037 7256 7348 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09036 7254 7350 7344 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09035 8144 7345 7254 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09034 7350 7351 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09033 8144 8063 7351 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09032 8144 7349 7348 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09031 7347 7350 7256 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09030 7255 7351 7347 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09029 8144 7346 7255 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09028 7346 7347 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09027 7344 7351 7346 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09026 8144 7344 7345 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09025 7345 7344 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09024 6260 6484 5976 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09023 5976 6480 6260 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09022 8144 6481 5976 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09021 7260 7358 7464 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09020 7259 7359 7260 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09019 8144 7357 7259 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09018 8144 3167 3168 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09017 3166 3168 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09016 8144 3165 3166 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09015 3260 3166 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09014 8144 3166 3260 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09013 8144 7458 7416 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09012 7416 7514 7507 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_09011 7734 7507 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_09010 508 509 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09009 503 510 506 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09008 8144 900 503 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09007 510 511 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09006 8144 1951 511 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_09005 8144 899 509 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09004 507 510 508 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09003 504 511 507 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09002 8144 505 504 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09001 505 507 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_09000 506 511 505 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08999 8144 506 900 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08998 900 506 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08997 7480 7725 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08996 8144 7724 7480 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08995 5836 5910 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08994 5835 5911 5836 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08993 8144 5909 5835 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08992 7731 7733 7698 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08991 8144 7956 7698 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08990 7698 7742 7731 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08989 7975 7731 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08988 6831 6830 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08987 6825 6833 6824 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08986 8144 6823 6825 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08985 6833 6832 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08984 8144 8063 6832 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08983 8144 6829 6830 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08982 6827 6833 6831 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08981 6828 6832 6827 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08980 8144 6826 6828 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08979 6826 6827 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08978 6824 6832 6826 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08977 8144 6824 6823 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08976 6823 6824 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08975 7901 7986 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08974 7899 7988 7980 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08973 8144 7979 7899 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08972 7988 7989 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08971 8144 8063 7989 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08970 8144 7985 7986 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08969 7984 7988 7901 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08968 7900 7989 7984 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08967 8144 7982 7900 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08966 7982 7984 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08965 7980 7989 7982 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08964 8144 7980 7979 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08963 7979 7980 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08962 8109 8067 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08961 8144 8068 8109 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08960 7268 7368 7471 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08959 7267 7369 7268 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08958 8144 7367 7267 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08957 6639 6652 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08956 8144 6636 6639 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08955 1813 4302 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08954 1813 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08953 8144 4575 1813 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08952 5166 5169 5058 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08951 8144 6850 5058 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08950 5058 5168 5166 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08949 5164 5166 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08948 1943 3348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08947 1943 2796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08946 8144 3542 1943 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08945 2339 2346 2279 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08944 8144 2616 2279 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08943 2279 2610 2339 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08942 2337 2339 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08941 6443 6564 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08940 6441 6565 6558 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08939 8144 6567 6441 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08938 6565 6566 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08937 8144 8063 6566 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08936 8144 6563 6564 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08935 6560 6565 6443 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08934 6442 6566 6560 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08933 8144 6559 6442 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08932 6559 6560 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08931 6558 6566 6559 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08930 8144 6558 6567 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08929 6567 6558 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08928 4539 4744 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08927 8144 4735 4539 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08926 4447 4539 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08925 6073 6071 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08924 8144 6070 6073 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08923 6332 6073 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08922 7301 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08921 7301 7398 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08920 8144 7884 7301 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08919 7114 7883 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08918 7114 7881 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08917 8144 7408 7114 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08916 6438 7559 6437 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08915 6437 7548 6534 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08914 6534 7550 6438 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08913 6438 6532 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08912 8144 6803 6438 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08911 6530 6534 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08910 3404 2718 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08909 3404 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08908 8144 4575 3404 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08907 2925 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08906 2925 2719 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08905 8144 4575 2925 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08904 7331 7332 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08903 8144 7330 7331 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08902 7737 7331 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08901 2152 3348 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08900 2152 3293 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08899 8144 3566 2152 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08898 8144 4511 3747 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08897 3747 4512 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08896 8144 3744 3747 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08895 3743 3747 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08894 8144 2870 2868 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08893 2870 3141 2748 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08892 2747 2872 2870 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08891 8144 3141 2872 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08890 2748 3348 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08889 8144 3315 2747 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08888 2868 2870 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08887 4508 4684 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08886 4505 4620 4680 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08885 8144 6549 4505 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08884 4620 4683 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08883 8144 8063 4683 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08882 8144 4681 4684 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08881 4619 4620 4508 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08880 4506 4683 4619 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08879 8144 4617 4506 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08878 4617 4619 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08877 4680 4683 4617 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08876 8144 4680 6549 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08875 6549 4680 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08874 7504 7747 7414 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08873 7414 7750 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08872 8144 7793 7504 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08871 7503 7504 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08870 5628 4548 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08869 5628 4707 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08868 8144 4529 5628 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08867 8144 4527 5628 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08866 7148 7147 6961 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_08865 6960 7305 7148 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_08864 8144 7301 6960 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_08863 6961 7158 8144 8144 pmos_3p3 L=0.28U W=4.77U AS=1.3356P AD=1.3356P PS=10.1U PD=10.1U 
Mtr_08862 7158 7891 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08861 7158 7892 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08860 8144 8187 7158 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08859 6956 7114 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08858 7108 7106 6956 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08857 8144 7104 7108 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08856 7885 7869 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08855 7885 7619 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08854 8144 8186 7885 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08853 5262 7149 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08852 5262 7887 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08851 8144 7130 5262 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08850 4024 5908 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08849 4024 3794 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08848 8144 4203 4024 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08847 3293 7528 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08846 3293 4173 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08845 8144 4172 3293 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08844 4007 6544 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08843 4007 6797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08842 8144 5648 4007 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08841 8144 5603 4007 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08840 7296 7869 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08839 7296 7398 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08838 8144 7892 7296 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08837 8048 3801 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08836 8048 3797 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08835 8144 7058 8048 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08834 8144 5908 8048 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08833 3033 4574 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08832 3033 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08831 8144 7356 3033 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08830 8144 6293 3033 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08829 8144 8059 8061 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08828 8144 8064 8065 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08827 8061 8065 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08826 8144 4498 4494 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08825 5092 4497 4412 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08824 4412 4498 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08823 4412 4494 5092 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08822 8144 4495 4412 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08821 4495 4497 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08820 4432 5417 4514 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_08819 4430 7787 4432 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_08818 4431 8048 4430 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_08817 8144 4429 4431 8144 pmos_3p3 L=0.28U W=3.09U AS=0.8652P AD=0.8652P PS=6.74U PD=6.74U 
Mtr_08816 4428 4514 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08815 5245 5868 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08814 5245 6172 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08813 8144 6921 5245 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08812 8144 7130 5245 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08811 4577 4572 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08810 4577 4575 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08809 8144 4573 4577 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08808 8144 4574 4577 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08807 7263 7970 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08806 8144 7957 7263 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08805 4957 6090 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08804 4956 6089 4957 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08803 8144 4955 4956 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08802 8144 5108 4676 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08801 4676 5938 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08800 8144 5606 4676 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08799 4921 4676 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08798 5834 7787 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08797 5913 5907 5834 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08796 8144 6801 5913 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08795 3222 3409 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08794 3410 4779 3222 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08793 8144 3857 3410 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08792 8051 8055 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08791 8144 8064 8051 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08790 2916 3379 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08789 8144 4540 2916 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08788 2918 2916 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08787 8144 3313 3309 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08786 4914 3310 3205 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08785 3205 3313 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08784 3205 3309 4914 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08783 8144 3311 3205 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08782 3311 3310 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08781 8144 8145 7868 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08780 7891 7868 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08779 8144 7868 7891 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08778 8144 7868 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08777 8144 7868 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08776 8144 8145 7864 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08775 7883 7864 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08774 8144 7864 7883 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08773 8144 7864 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08772 8144 7864 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08771 8144 8145 8146 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08770 8184 8146 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08769 8144 8146 8184 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08768 8144 8146 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08767 8144 8146 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08766 8144 8145 7870 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08765 7869 7870 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08764 8144 7870 7869 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08763 8144 7870 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08762 8144 7870 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08761 8144 5680 5681 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08760 8145 5681 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08759 8144 5681 8145 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08758 8144 5681 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08757 8144 5681 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08756 8144 3405 3406 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08755 3406 4276 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08754 8144 3404 3406 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08753 3641 3406 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08752 8144 3857 2780 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08751 2780 2943 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08750 3177 4575 2780 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08749 2779 2937 3177 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08748 2780 2938 2779 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08747 564 1372 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08746 8144 1157 564 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08745 565 564 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08744 1959 1957 1845 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08743 1845 1956 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08742 8144 1962 1959 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08741 2167 1959 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08740 8144 969 573 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08739 5483 573 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08738 8144 573 5483 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08737 8144 573 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08736 8144 573 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08735 8144 969 970 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08734 5942 970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08733 8144 970 5942 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08732 8144 970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08731 8144 970 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08730 8144 579 578 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08729 969 578 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08728 8144 578 969 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08727 8144 578 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08726 8144 578 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08725 8144 384 382 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08724 5654 382 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08723 8144 382 5654 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08722 8144 382 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08721 8144 382 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08720 8144 384 383 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08719 5447 383 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08718 8144 383 5447 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08717 8144 383 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08716 8144 383 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08715 8144 386 385 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08714 384 385 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08713 8144 385 384 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08712 8144 385 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08711 8144 385 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08710 8144 6312 6313 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08709 7352 6313 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08708 8144 6313 7352 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08707 8144 6313 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08706 8144 6313 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08705 8144 6312 6306 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08704 7041 6306 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08703 8144 6306 7041 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08702 8144 6306 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08701 8144 6306 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08700 8144 5916 5915 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08699 6312 5915 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08698 8144 5915 6312 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08697 8144 5915 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08696 8144 5915 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08695 5442 5633 5441 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08694 5441 5444 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08693 8144 7068 5442 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08692 5440 5442 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08691 8144 7058 3605 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08690 3605 3801 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08689 8144 5908 3605 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08688 5633 3605 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08687 8144 1375 1376 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08686 1376 1377 1590 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08685 8144 5509 5039 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08684 5039 5037 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08683 8144 5038 5039 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08682 5036 5039 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08681 8144 1583 1579 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08680 1579 2022 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08679 8144 1576 1579 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08678 3156 1579 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08677 8144 4193 4196 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08676 4196 4192 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08675 8144 4438 4196 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08674 4191 4196 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08673 8144 6076 2883 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08672 8144 8064 2884 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08671 2883 2884 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08670 8144 4663 4659 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08669 4662 4658 4587 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08668 4587 4663 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08667 4587 4659 4662 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08666 8144 4660 4587 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08665 4660 4658 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08664 8144 4068 959 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08663 959 6311 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08662 959 4572 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08661 8144 3857 959 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08660 1375 959 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08659 930 932 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08658 926 933 927 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08657 8144 1113 926 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08656 933 934 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08655 8144 3834 934 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08654 8144 935 932 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08653 931 933 930 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08652 928 934 931 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08651 8144 929 928 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08650 929 931 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08649 927 934 929 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08648 8144 927 1113 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08647 1113 927 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08646 5853 6127 5854 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08645 5852 6145 5853 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08644 8144 6618 5852 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08643 7790 7788 7792 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08642 7792 7791 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08641 8144 8040 7790 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08640 7789 7790 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08639 8144 4068 1186 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08638 1186 4295 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08637 1186 5648 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08636 8144 4067 1186 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08635 1390 1186 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08634 8144 1618 1442 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08633 1442 1617 1619 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08632 3224 3650 3268 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08631 3223 3664 3224 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08630 8144 3267 3223 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08629 4554 4754 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08628 4550 4634 4752 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08627 8144 4760 4550 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08626 4634 4755 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08625 8144 5864 4755 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08624 8144 4759 4754 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08623 4633 4634 4554 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08622 4551 4755 4633 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08621 8144 4631 4551 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08620 4631 4633 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08619 4752 4755 4631 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08618 8144 4752 4760 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08617 4760 4752 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08616 4600 4734 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08615 4735 6363 4600 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08614 8144 6359 4735 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08613 4244 4449 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08612 8144 4448 4244 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08611 6156 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08610 8144 6396 6156 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08609 6158 7633 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08608 8144 6652 6158 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08607 7819 7820 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08606 7815 7822 7814 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08605 8144 8071 7815 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08604 7822 7823 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08603 8144 7821 7823 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08602 8144 8070 7820 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08601 7818 7822 7819 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08600 7816 7823 7818 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08599 8144 7817 7816 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08598 7817 7818 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08597 7814 7823 7817 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08596 8144 7814 8071 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08595 8071 7814 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08594 7420 7797 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08593 7523 7798 7420 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08592 8144 8139 7523 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08591 5160 5435 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08590 5160 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08589 8144 7352 5160 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08588 4448 4749 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08587 8144 4955 4448 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08586 6615 8179 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08585 8144 7872 6615 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08584 5148 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08583 5148 1565 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08582 8144 6609 5148 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08581 4518 4306 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08580 4518 1565 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08579 8144 6802 4518 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08578 8144 2710 2715 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08577 2713 2712 2957 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08576 2714 2942 2713 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08575 2715 2932 2714 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08574 342 3622 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08573 8144 1150 342 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08572 159 365 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08571 8144 166 159 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08570 8144 3147 3315 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08569 3147 3780 3068 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08568 3069 3070 3147 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08567 8144 3780 3070 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08566 3068 3353 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08565 8144 3602 3069 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08564 3315 3147 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08563 8144 3359 4510 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08562 3359 3780 3217 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08561 3216 3363 3359 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08560 8144 3780 3363 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08559 3217 3361 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08558 8144 5180 3216 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08557 4510 3359 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08556 8144 3350 3348 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08555 3350 3780 3214 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08554 3213 3355 3350 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08553 8144 3780 3355 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08552 3214 3353 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08551 8144 4030 3213 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08550 3348 3350 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08549 5562 5563 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08548 5562 7361 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08547 8144 7041 5562 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08546 5495 5498 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08545 8144 5706 5495 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08544 1543 6796 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08543 1543 4068 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08542 8144 6609 1543 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08541 1469 5099 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08540 8144 1466 1469 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08539 1467 1469 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08538 2600 3553 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08537 8144 2798 2600 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08536 2599 2600 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08535 3547 3562 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08534 3549 3757 3544 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08533 3544 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08532 8144 3545 3550 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08531 3550 3546 3548 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08530 3548 3547 3549 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08529 3549 3562 3551 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08528 3551 4426 3550 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08527 8144 3556 3545 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08526 3986 3549 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08525 3560 3562 8144 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08524 3563 3995 3557 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08523 3557 3556 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08522 8144 3558 3564 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08521 3564 3559 3561 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08520 3561 3560 3563 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08519 3563 3562 3565 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08518 3565 3754 3564 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08517 8144 3556 3558 8144 pmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08516 4141 3563 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08515 7904 7996 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08514 7902 7997 7991 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08513 8144 8000 7902 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08512 7997 7998 8144 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08511 8144 8063 7998 8144 pmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08510 8144 7999 7996 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08509 7995 7997 7904 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08508 7903 7998 7995 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08507 8144 7992 7903 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08506 7992 7995 8144 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08505 7991 7998 7992 8144 pmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08504 8144 7991 8000 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08503 8000 7991 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08502 5418 5417 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08501 6784 5432 5418 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08500 8144 5416 6784 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08499 2219 2227 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08498 8144 4518 2219 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08497 2437 2219 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08496 7401 7639 7303 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08495 7303 8180 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08494 8144 7633 7401 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08493 7302 7401 8144 8144 pmos_3p3 L=0.28U W=3.19U AS=0.8932P AD=0.8932P PS=6.95U PD=6.95U 
Mtr_08492 8144 6573 6843 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08491 6573 6867 6447 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08490 6446 6575 6573 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08489 8144 6867 6575 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08488 6447 6663 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08487 8144 6838 6446 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08486 6843 6573 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08485 8144 6866 6863 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08484 6866 6867 6868 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08483 6865 6869 6866 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08482 8144 6867 6869 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08481 6868 7283 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08480 8144 6864 6865 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08479 6863 6866 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08478 8144 6605 6600 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08477 6605 6867 6455 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08476 6454 6606 6605 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08475 8144 6867 6606 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08474 6455 6632 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08473 8144 6602 6454 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08472 6600 6605 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08471 8144 179 177 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08470 179 4538 180 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08469 178 181 179 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08468 8144 4538 181 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08467 180 187 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08466 8144 4540 178 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08465 177 179 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08464 8144 6902 6900 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08463 6902 7867 6903 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08462 6901 6904 6902 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08461 8144 7867 6904 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08460 6903 6988 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08459 8144 7119 6901 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08458 6900 6902 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08457 8144 7387 7893 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08456 7387 7867 7290 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08455 7291 7292 7387 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08454 8144 7867 7292 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08453 7290 7777 8144 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08452 8144 7604 7291 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08451 7893 7387 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08450 4517 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08449 4517 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08448 8144 5648 4517 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08447 5147 7051 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08446 5147 4310 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08445 8144 5483 5147 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08444 6791 6794 8144 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08443 8144 7343 6791 8144 pmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08442 7007 6791 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08441 1932 2152 1839 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08440 1839 2608 1932 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08439 8144 2616 1839 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08438 2617 2827 2618 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08437 8144 2616 2618 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08436 2618 3307 2617 8144 pmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08435 2816 2617 8144 8144 pmos_3p3 L=0.28U W=4.03U AS=1.1284P AD=1.1284P PS=8.63U PD=8.63U 
Mtr_08434 7228 7333 7229 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08433 7229 7336 7335 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08432 8185 7334 7228 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08431 7520 7335 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08430 660 923 662 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08429 8185 662 659 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08428 8185 923 663 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08427 661 3537 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08426 662 663 661 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08425 8185 676 660 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08424 659 662 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08423 257 923 258 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08422 8185 258 256 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08421 8185 923 260 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08420 259 3532 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08419 258 260 259 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08418 8185 266 257 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08417 256 258 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08416 3376 4293 3377 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08415 3377 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08414 3378 5648 3376 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08413 6728 7867 6896 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08412 8185 6896 6893 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08411 8185 7867 6898 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08410 6729 7061 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08409 6896 6898 6729 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08408 8185 7112 6728 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08407 6893 6896 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08406 7116 7867 7117 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08405 8185 7117 7408 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08404 8185 7867 7120 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08403 7118 7349 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08402 7117 7120 7118 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08401 8185 7379 7116 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_08400 7408 7117 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08399 1585 5654 1584 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08398 1584 4295 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08397 1582 5942 1585 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08396 1583 7051 1582 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08395 1197 1710 1198 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08394 1198 1455 1291 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08393 8185 1729 1197 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08392 1293 1291 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08391 3718 3722 3719 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08390 3719 3717 3718 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08389 8185 3971 3719 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08388 8185 7147 6651 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08387 6651 7140 6650 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08386 6648 6650 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08385 6124 6907 6123 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08384 6123 7361 6124 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08383 8185 6576 6123 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08382 6133 6124 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08381 8185 7872 7684 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08380 7684 8179 7873 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08379 7874 7873 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08378 3977 4009 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08377 8185 7787 3977 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08376 3977 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08375 8185 8045 3977 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08374 3972 3977 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08373 2825 4574 2826 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08372 2826 6797 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08371 2823 7353 2825 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08370 2822 2824 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_08369 2824 6484 2823 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08368 8185 5139 5141 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08367 5141 5440 5142 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08366 5140 5142 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08365 1 62 4644 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08364 8185 1928 1 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08363 2 1284 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08362 4644 61 2 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08361 8185 1284 62 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08360 61 1928 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08359 7483 7723 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08358 7482 7480 7483 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08357 8185 7481 7482 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08356 7492 7482 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08355 8185 5942 2446 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08354 2446 7356 2445 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08353 2894 2445 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08352 8185 5654 815 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08351 815 6609 941 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08350 1352 941 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08349 4692 6821 4691 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08348 4691 5406 4692 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08347 8185 6809 4691 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08346 4690 4692 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08345 762 562 434 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08344 434 764 762 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08343 8185 1364 434 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08342 4741 4737 4740 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08341 4740 4738 4741 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08340 8185 4739 4740 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08339 4983 4741 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08338 5697 6156 5699 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08337 5699 6157 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08336 5698 6166 5697 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08335 5695 5696 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_08334 5696 7880 5698 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08333 5154 8047 5155 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08332 5155 5907 5154 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08331 8185 6541 5155 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08330 8185 3033 2949 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08329 2949 4470 2948 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08328 2947 2948 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08327 4830 7026 4831 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08326 4831 6797 4930 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08325 8185 6544 4830 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08324 5907 4930 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08323 8185 7883 5741 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08322 5741 7408 5742 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08321 5740 5742 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08320 3053 3405 3054 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08319 3054 3177 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08318 3052 4276 3053 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08317 3872 3178 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_08316 3178 3404 3052 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08315 2007 4574 2009 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08314 2009 4068 2008 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08313 8185 2492 2007 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08312 2006 2008 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08311 49 558 50 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08310 50 559 167 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08309 8185 1362 49 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08308 166 167 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08307 4351 4535 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08306 4350 4532 4534 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08305 4349 4536 4531 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08304 8185 4720 4349 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08303 8185 5864 4536 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08302 4532 4536 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08301 8185 4721 4535 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08300 4534 4536 4351 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08299 4533 4534 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08298 8185 4533 4350 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08297 4531 4532 4533 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08296 4720 4531 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08295 8185 4531 4720 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08294 5625 7356 5627 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08293 5627 6802 5626 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08292 8185 5624 5625 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08291 7798 5626 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08290 1161 1996 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08289 8185 2698 1161 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08288 1161 1891 1588 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08287 1588 2926 1161 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08286 6237 6907 6238 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08285 6238 7398 6397 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08284 8185 7891 6237 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08283 6396 6397 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08282 2118 5654 2117 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08281 2117 4293 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08280 2116 5483 2118 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08279 2256 2257 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_08278 2257 3857 2116 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08277 3256 4051 3257 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08276 3257 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08275 3255 7026 3256 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08274 3635 3397 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_08273 3397 5624 3255 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08272 2330 2601 2331 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08271 2331 2344 2330 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08270 8185 2589 2331 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08269 2596 2330 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08268 8185 6152 5904 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08267 5832 5904 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08266 8185 5904 5832 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08265 8185 5904 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08264 8144 5904 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08263 8185 5961 5903 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08262 5831 5903 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08261 8185 5903 5831 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08260 8185 5903 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08259 8144 5903 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08258 8185 6152 2021 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08257 3834 2021 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08256 8185 2021 3834 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08255 8185 2021 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08254 8144 2021 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08253 8185 6152 2020 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08252 2019 2020 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08251 8185 2020 2019 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08250 8185 2020 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08249 8144 2020 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08248 8185 6152 1810 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08247 1809 1810 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08246 8185 1810 1809 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08245 8185 1810 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08244 8144 1810 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08243 8185 5961 1808 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08242 1807 1808 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08241 8185 1808 1807 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08240 8185 1808 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08239 8144 1808 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08238 8185 6152 1953 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08237 3708 1953 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08236 8185 1953 3708 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08235 8185 1953 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08234 8144 1953 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08233 8185 6152 1952 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08232 1951 1952 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08231 8185 1952 1951 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08230 8185 1952 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08229 8144 1952 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08228 8185 6152 1748 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08227 1772 1748 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08226 8185 1748 1772 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08225 8185 1748 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08224 8144 1748 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08223 8185 5961 1747 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08222 1746 1747 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08221 8185 1747 1746 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08220 8185 1747 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08219 8144 1747 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08218 6181 7151 6180 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08217 6179 6672 6181 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08216 6180 6658 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08215 6177 6181 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08214 8185 6668 6179 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08213 6179 6178 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08212 8185 190 189 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08211 57 189 188 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08210 8185 1699 57 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08209 187 188 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08208 8185 188 187 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08207 3182 2039 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08206 8185 2041 3182 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08205 395 483 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08204 394 484 480 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08203 393 485 478 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08202 8185 676 393 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08201 8185 1951 485 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08200 484 485 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08199 8185 659 483 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08198 480 485 395 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08197 479 480 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08196 8185 479 394 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08195 478 484 479 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08194 676 478 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08193 8185 478 676 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08192 6997 7000 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08191 6996 6999 6998 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08190 6993 7001 6994 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08189 8185 6992 6993 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08188 8185 8063 7001 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08187 6999 7001 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08186 8185 7777 7000 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08185 6998 7001 6997 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08184 6995 6998 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08183 8185 6995 6996 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08182 6994 6999 6995 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08181 6992 6994 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08180 8185 6994 6992 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08179 1475 3969 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08178 1474 1473 1475 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08177 1107 1115 1109 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08176 1109 1114 1108 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08175 1108 1113 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08174 1106 1111 1109 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08173 8185 1110 1106 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08172 8185 1116 1107 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08171 1325 1109 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08170 7965 7490 7491 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08169 7491 7497 7965 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08168 8185 7489 7491 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08167 2349 4172 2350 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08166 2350 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08165 2796 7549 2349 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08164 7081 7084 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08163 7083 7085 7082 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08162 7078 7086 7079 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08161 8185 7272 7078 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08160 8185 7821 7086 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08159 7085 7086 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08158 8185 7271 7084 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08157 7082 7086 7081 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08156 7080 7082 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08155 8185 7080 7083 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08154 7079 7085 7080 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08153 7272 7079 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08152 8185 7079 7272 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08151 7781 7779 7663 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08150 7663 7778 7781 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08149 8185 7777 7663 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08148 8052 7781 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08147 7465 7464 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08146 8136 7765 7465 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08145 3059 3186 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08144 3267 3187 3059 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08143 8185 1157 1159 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_08142 1159 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_08141 2022 1158 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08140 1159 2227 1158 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_08139 1158 2926 1159 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_08138 4953 6090 4839 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08137 4839 6089 4953 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08136 8185 6341 4839 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08135 7972 7977 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08134 7974 7976 7973 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08133 7968 7978 7969 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08132 8185 8008 7968 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08131 8185 8063 7978 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08130 7976 7978 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08129 8185 7975 7977 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08128 7973 7978 7972 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08127 7971 7973 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08126 8185 7971 7974 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08125 7969 7976 7971 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08124 8008 7969 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08123 8185 7969 8008 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08122 5363 5508 5362 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08121 5362 5507 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08120 5361 5503 5363 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08119 5504 7880 5361 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08118 7109 7408 7111 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08117 7111 7892 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08116 7110 7883 7109 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08115 828 2719 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08114 957 7051 828 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08113 1902 1589 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08112 8185 1587 1902 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08111 1902 1892 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08110 8185 1588 1902 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08109 1816 1617 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08108 8185 1618 1816 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08107 1816 1615 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08106 8185 1616 1816 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08105 8185 3553 2990 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08104 2990 3543 3103 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08103 3102 3103 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08102 6223 6321 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08101 6222 6322 6317 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08100 6221 6323 6314 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08099 8185 6344 6221 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08098 8185 8063 6323 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08097 6322 6323 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08096 8185 6319 6321 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08095 6317 6323 6223 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08094 6316 6317 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08093 8185 6316 6222 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08092 6314 6322 6316 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08091 6344 6314 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08090 8185 6314 6344 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08089 2545 2669 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08088 2546 2670 2667 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08087 2544 2671 2663 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08086 8185 6076 2544 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08085 8185 3708 2671 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08084 2670 2671 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_08083 8185 2668 2669 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_08082 2667 2671 2545 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08081 2664 2667 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08080 8185 2664 2546 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08079 2663 2670 2664 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08078 6076 2663 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08077 8185 2663 6076 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08076 6053 6051 6052 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08075 6052 6778 6053 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08074 8185 7314 6052 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08073 6050 6053 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08072 8185 5426 5306 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08071 5306 5629 5427 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08070 5618 5427 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08069 5639 5637 5640 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08068 5638 5642 5639 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08067 5640 5644 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08066 6095 5639 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08065 8185 5653 5638 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08064 5638 5641 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_08063 5367 6636 5368 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08062 5368 6909 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08061 5366 6921 5367 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08060 5508 7130 5366 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08059 5355 6921 5354 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08058 5354 7880 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08057 6629 7130 5355 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08056 7472 7471 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08055 8156 7566 7472 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_08054 7632 7893 7631 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08053 7631 7630 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08052 7876 8184 7632 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08051 3044 3579 3045 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08050 3045 3356 3138 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08049 8185 3582 3044 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08048 3137 3138 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_08047 1201 1710 1200 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08046 1200 1455 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08045 1295 1729 1201 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08044 8185 1301 1205 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08043 1205 5395 1299 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08042 1719 1299 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08041 3756 4511 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08040 3755 4512 3756 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08039 8185 4510 3755 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08038 3754 3755 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08037 3332 3763 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08036 3331 4424 3332 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08035 8185 4510 3331 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08034 3330 3331 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08033 5028 6177 4862 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08032 4862 5504 5028 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08031 8185 5026 4862 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08030 5027 5028 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08029 5252 6654 5251 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08028 5251 8179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08027 5250 7633 5252 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08026 5249 7130 5250 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08025 5692 6154 5694 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08024 5694 5865 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08023 5693 6158 5692 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08022 6241 6647 6242 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08021 6242 6906 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08020 6403 6632 6241 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08019 2104 2239 2105 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08018 2105 2238 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08017 2467 3172 2104 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08016 8185 7880 5356 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08015 5356 5503 5499 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08014 5500 5499 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08013 6733 7881 6734 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08012 6734 7398 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08011 6905 8184 6733 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08010 4673 4670 4672 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08009 8185 7029 4673 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08008 4674 4900 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08007 4672 4671 4674 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08006 8185 4900 4670 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08005 4671 7029 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08004 8185 4078 3653 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08003 8185 3651 3653 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08002 3653 3851 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_08001 3650 3653 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_08000 8185 3073 3194 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07999 3194 3650 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07998 3197 3194 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07997 8185 7885 7692 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07996 7692 7889 7886 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07995 8171 7886 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07994 6168 6652 6170 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07993 6170 7121 6169 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07992 8185 6636 6168 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07991 6378 6169 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07990 7516 7761 7515 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07989 7515 7760 7516 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07988 8185 8008 7515 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07987 7514 7516 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07986 3457 3578 4502 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07985 8185 3575 3457 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07984 3456 3577 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07983 4502 3574 3456 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07982 8185 3577 3578 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07981 3574 3575 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07980 8185 3175 2921 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07979 7353 2921 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07978 8185 2921 7353 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07977 8185 2921 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07976 8144 2921 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07975 8185 3175 781 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07974 7051 781 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07973 8185 781 7051 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07972 8185 781 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07971 8144 781 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07970 8185 3175 3176 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07969 6293 3176 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07968 8185 3176 6293 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07967 8185 3176 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07966 8144 3176 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07965 8185 3175 2457 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07964 6796 2457 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07963 8185 2457 6796 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07962 8185 2457 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07961 8144 2457 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07960 8185 3175 3169 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07959 6544 3169 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07958 8185 3169 6544 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07957 8185 3169 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07956 8144 3169 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07955 8185 369 368 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07954 3175 368 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07953 8185 368 3175 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07952 8185 368 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07951 8144 368 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07950 3051 3844 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07949 3172 4295 3051 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07948 3050 3399 3172 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07947 8185 3170 3050 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07946 3050 3171 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07945 8185 4292 3869 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07944 3869 3867 3870 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07943 3868 3870 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07942 8185 1184 1183 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07941 3857 1183 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07940 8185 1183 3857 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07939 8185 1183 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07938 8144 1183 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07937 8185 1184 1185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07936 4075 1185 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07935 8185 1185 4075 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07934 8185 1185 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07933 8144 1185 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07932 8185 963 964 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07931 1184 964 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07930 8185 964 1184 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07929 8185 964 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07928 8144 964 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07927 6779 6775 6683 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07926 8185 7500 6777 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07925 6683 6777 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07924 41 553 40 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07923 40 365 160 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07922 8185 166 41 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07921 334 160 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07920 2074 7026 2075 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07919 2075 6543 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07918 2073 7353 2074 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07917 2198 2197 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07916 2197 6080 2073 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07915 2897 2896 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07914 7058 4067 2897 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07913 2895 6796 7058 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07912 8185 2898 2895 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07911 2895 2894 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07910 2486 2484 2488 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07909 2488 2485 2487 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07908 8185 2947 2486 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07907 2955 2487 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07906 4686 7029 4687 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07905 4687 5406 4686 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07904 8185 6798 4687 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07903 4685 4686 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07902 5778 5949 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07901 5779 5950 5948 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07900 5777 5951 5946 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07899 8185 6375 5777 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07898 8185 7821 5951 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07897 5950 5951 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07896 8185 6374 5949 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07895 5948 5951 5778 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07894 5947 5948 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07893 8185 5947 5779 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07892 5946 5950 5947 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07891 6375 5946 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07890 8185 5946 6375 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07889 5226 5238 5225 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07888 5225 6629 5226 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07887 8185 5223 5225 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07886 4656 4654 4663 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07885 8185 6524 4656 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07884 4657 4895 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07883 4663 4655 4657 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07882 8185 4895 4654 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07881 4655 6524 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07880 1266 7026 1268 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07879 1268 6543 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07878 1267 5624 1266 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07877 1593 1380 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07876 1380 3857 1267 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07875 1182 4068 1181 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07874 1181 6802 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07873 1180 4306 1182 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07872 2252 1179 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07871 1179 3857 1180 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07870 3461 3783 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07869 3586 3782 3461 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07868 3342 3780 3343 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07867 3341 3579 3342 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07866 3343 4255 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07865 3340 3342 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07864 8185 3587 3341 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07863 3341 3774 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07862 301 304 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07861 300 303 302 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07860 297 305 298 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07859 8185 709 297 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07858 8185 1772 305 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07857 303 305 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07856 8185 710 304 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07855 302 305 301 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07854 299 302 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07853 8185 299 300 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07852 298 303 299 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07851 709 298 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07850 8185 298 709 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07849 5192 5193 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07848 5190 5195 5191 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07847 5187 5194 5186 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07846 8185 5197 5187 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07845 8185 5864 5194 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07844 5195 5194 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07843 8185 5196 5193 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07842 5191 5194 5192 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07841 5189 5191 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07840 8185 5189 5190 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07839 5186 5195 5189 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07838 5197 5186 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07837 8185 5186 5197 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07836 5438 7059 5313 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07835 5313 6294 5438 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07834 8185 5437 5313 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07833 5436 5438 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07832 6016 6520 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07831 6015 6618 6016 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07830 6031 6383 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07829 6614 6145 6031 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07828 4580 4583 4382 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07827 4382 5037 4580 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07826 8185 4579 4382 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07825 4474 4580 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07824 4315 4583 4316 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07823 4316 5041 4315 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07822 8185 4317 4316 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07821 3266 3419 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07820 3423 3264 3266 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07819 3781 3780 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07818 3782 4543 3781 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07817 2057 5401 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07816 2813 2159 2057 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07815 3122 3123 2997 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07814 2997 3569 3122 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07813 8185 3567 2997 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07812 3121 3122 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07811 5803 7872 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07810 5866 6396 5803 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07809 5341 6383 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07808 5489 5485 5341 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07807 5346 6654 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07806 5494 6396 5346 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07805 4852 6383 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07804 5486 5202 4852 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07803 5739 7887 5738 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07802 5738 5879 5739 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07801 8185 5878 5738 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07800 5737 5739 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07799 3504 3871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07798 3664 3665 3504 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07797 3060 3268 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07796 3264 3192 3060 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07795 443 1150 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07794 553 6363 443 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07793 5754 7752 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07792 5902 6285 5754 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07791 5753 6286 5902 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07790 8185 5898 5753 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07789 5752 6549 5902 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07788 8185 6284 5752 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07787 6 1924 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07786 1929 1711 6 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07785 7676 7834 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07784 7675 7832 7831 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07783 7674 7833 7826 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07782 8185 7824 7674 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07781 8185 8166 7833 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07780 7832 7833 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07779 8185 7829 7834 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07778 7831 7833 7676 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07777 7827 7831 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07776 8185 7827 7675 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07775 7826 7832 7827 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07774 7824 7826 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07773 8185 7826 7824 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07772 5284 7352 5285 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07771 5285 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07770 5388 5387 5284 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07769 8185 955 761 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07768 8185 956 761 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07767 761 762 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07766 943 761 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07765 8054 7029 7030 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07764 7030 7058 8054 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07763 8185 7048 7030 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07762 1251 4573 1250 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07761 1250 6311 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07760 1559 4067 1251 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07759 5807 7884 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07758 5868 8184 5807 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07757 4288 4583 4289 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07756 4289 5031 4288 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07755 8185 4286 4289 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07754 4287 4288 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07753 8185 7323 7170 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07752 7170 7325 7324 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07751 7319 7324 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07750 8185 4007 3002 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07749 3002 3146 3140 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07748 3139 3140 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07747 8017 8016 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07746 8013 8018 8014 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07745 8011 8019 8010 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07744 8185 8021 8011 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07743 8185 8063 8019 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07742 8018 8019 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07741 8185 8020 8016 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07740 8014 8019 8017 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07739 8012 8014 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07738 8185 8012 8013 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07737 8010 8018 8012 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07736 8021 8010 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07735 8185 8010 8021 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07734 8185 6359 5328 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07733 5455 8122 5325 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07732 5452 5665 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_07731 5325 5450 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07730 8185 6359 5450 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_07729 5449 5455 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_07728 5328 5658 5327 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07727 5327 5665 5455 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07726 5455 5452 5326 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07725 5326 5453 5328 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07724 399 923 495 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07723 8185 495 496 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07722 8185 923 453 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07721 400 3978 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07720 495 453 400 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07719 8185 497 399 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07718 496 495 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07717 731 923 921 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07716 8185 921 920 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07715 8185 923 925 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07714 734 4012 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07713 921 925 734 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07712 8185 1111 731 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07711 920 921 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07710 699 923 698 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07709 8185 698 697 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07708 8185 923 701 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07707 700 4160 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07706 698 701 700 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07705 8185 703 699 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07704 697 698 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07703 726 923 728 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07702 8185 728 724 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07701 8185 923 727 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07700 729 4176 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07699 728 727 729 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07698 8185 725 726 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07697 724 728 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07696 288 923 290 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07695 8185 290 287 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07694 8185 923 291 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07693 289 3999 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07692 290 291 289 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07691 8185 512 288 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07690 287 290 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07689 2892 4573 2893 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07688 2893 6311 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07687 5168 4293 2892 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07686 1254 2013 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07685 1368 3148 1254 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07684 6690 6797 6691 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07683 6691 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07682 6689 6796 6690 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07681 7328 6792 6689 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07680 8185 3229 2059 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07679 2059 2166 2165 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07678 2355 2165 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07677 7252 7797 7177 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07676 7177 7798 7252 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07675 8185 7777 7177 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07674 5309 5629 5310 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07673 5310 5628 5433 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07672 8185 5434 5309 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07671 5432 5433 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07670 308 923 307 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07669 8185 307 306 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07668 8185 923 310 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07667 309 2402 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07666 307 310 309 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07665 8185 529 308 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07664 306 307 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07663 687 1332 892 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07662 8185 892 890 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07661 8185 1332 894 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07660 690 3537 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07659 892 894 690 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07658 8185 1048 687 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07657 890 892 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07656 1040 1332 1039 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07655 8185 1039 1038 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07654 8185 1332 1042 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07653 1041 3532 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07652 1039 1042 1041 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07651 8185 1043 1040 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07650 1038 1039 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07649 682 1332 887 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07648 8185 887 885 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07647 8185 1332 889 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07646 683 3978 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07645 887 889 683 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07644 8185 1304 682 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07643 885 887 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07642 5098 5108 5097 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07641 5097 6801 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07640 5096 5938 5098 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07639 5110 5606 5096 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07638 3025 4167 3024 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07637 3024 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07636 3379 5624 3025 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07635 6190 6667 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07634 8185 6188 6190 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07633 6190 7299 6191 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07632 6191 6189 6190 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07631 8185 2941 2244 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07630 8185 2242 2244 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07629 2244 2241 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07628 3656 2244 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07627 3806 5447 3807 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07626 3807 4167 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07625 3805 7051 3806 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07624 3804 5664 3805 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07623 2810 4172 2812 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07622 2812 4173 2811 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07621 8185 7528 2810 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07620 2809 2811 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07619 1922 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07618 1924 2602 1922 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07617 1923 2141 1924 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07616 8185 3737 1923 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07615 1923 2136 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07614 1665 6359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07613 8185 2698 1665 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07612 1665 1887 1893 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07611 1893 2926 1665 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07610 6701 7500 7061 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07609 8185 7500 6808 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07608 6702 7345 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07607 7061 6808 6702 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07606 8185 6804 6701 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07605 8185 2941 2945 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07604 8185 2946 2945 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07603 2945 2942 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07602 3645 2945 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07601 8185 3556 2368 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07600 2370 3562 2363 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07599 2367 2379 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_07598 2363 2364 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07597 8185 3556 2364 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_07596 2635 2370 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_07595 2368 2365 2366 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07594 2366 2379 2370 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07593 2370 2367 2369 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07592 2369 2843 2368 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07591 8185 3556 2360 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07590 2358 2352 2354 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07589 2357 2379 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_07588 2354 2353 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07587 8185 3556 2353 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_07586 3108 2358 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_07585 2360 2355 2356 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07584 2356 2379 2358 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07583 2358 2357 2359 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07582 2359 2840 2360 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_07581 8185 4197 4199 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07580 8047 4199 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07579 8185 4199 8047 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07578 8185 4199 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07577 8144 4199 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07576 8185 3771 3772 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07575 4197 3772 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07574 8185 3772 4197 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07573 8185 3772 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07572 8144 3772 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07571 5651 5654 5652 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07570 5652 5648 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07569 5649 6796 5651 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07568 5929 5650 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07567 5650 6375 5649 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07566 6486 7500 7280 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07565 8185 7500 6488 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07564 6487 6974 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07563 7280 6488 6487 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07562 8185 6485 6486 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07561 8188 8186 8189 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07560 8189 8187 8188 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07559 8185 8184 8189 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07558 366 3391 367 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07557 367 1150 366 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07556 8185 3393 367 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07555 365 366 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07554 8185 5917 5756 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07553 5756 5902 5901 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07552 5830 5901 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07551 8185 1346 1231 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07550 1231 1348 1347 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07549 4025 1347 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07548 8185 4197 4008 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07547 7787 4008 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07546 8185 4008 7787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07545 8185 4008 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07544 8144 4008 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07543 5104 5105 5121 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07542 8185 5938 5104 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07541 5103 5108 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07540 5121 5102 5103 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07539 8185 5108 5105 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07538 5102 5938 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07537 5884 6270 5792 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07536 5791 7550 5884 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07535 5792 6271 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07534 5817 5884 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07533 8185 7548 5791 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07532 5791 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07531 402 1115 501 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07530 501 1114 403 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07529 403 685 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07528 401 497 501 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07527 8185 1110 401 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07526 8185 498 402 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07525 1738 501 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07524 6810 7061 6703 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07523 6703 6835 6810 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07522 8185 7053 6703 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07521 6809 6810 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07520 2526 2631 2633 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07519 2633 2836 2527 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07518 2527 3744 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07517 2525 2636 2633 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07516 8185 3112 2525 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07515 8185 2630 2526 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07514 2830 2633 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07513 1193 1286 1284 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07512 8185 2132 1193 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07511 1194 2133 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07510 1284 1283 1194 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07509 8185 2133 1286 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07508 1283 2132 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07507 8185 4951 4711 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07506 7343 4711 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07505 8185 4711 7343 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07504 8185 4711 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07503 8144 4711 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07502 8185 4951 4952 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07501 5574 4952 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07500 8185 4952 5574 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07499 8185 4952 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07498 8144 4952 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07497 8185 4525 4526 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07496 4951 4526 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07495 8185 4526 4951 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07494 8185 4526 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07493 8144 4526 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07492 5801 6156 5802 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07491 5802 6403 5964 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07490 8185 6166 5801 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07489 5865 5964 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07488 8185 7891 7202 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07487 7202 7398 7377 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07486 7283 7377 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07485 2606 2809 2511 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07484 2511 3320 2606 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07483 8185 3315 2511 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07482 2605 2606 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07481 3555 3552 3445 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07480 3445 3748 3555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07479 8185 3553 3445 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07478 3740 3555 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07477 3810 3812 3811 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07476 3811 3809 3810 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07475 8185 7314 3811 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07474 4737 3810 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07473 7767 6524 6525 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07472 6525 7058 7767 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07471 8185 7012 6525 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07470 5374 5373 5277 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07469 5276 7550 5374 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07468 5277 5551 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07467 5372 5374 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07466 8185 7548 5276 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07465 5276 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_07464 1367 1571 1252 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07463 1252 1570 1367 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07462 8185 1364 1252 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07461 1365 1367 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07460 576 5940 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07459 8185 2262 576 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07458 3742 3743 3741 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07457 3741 3740 3742 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07456 8185 4141 3741 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07455 4157 3742 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07454 1755 2178 1650 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07453 1650 2179 1755 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07452 8185 1962 1650 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07451 2170 1755 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07450 3289 3720 3288 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07449 3288 4492 3289 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07448 8185 3286 3288 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07447 3287 3289 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07446 315 318 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07445 314 317 316 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07444 311 319 312 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07443 8185 725 311 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07442 8185 1772 319 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07441 317 319 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07440 8185 724 318 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07439 316 319 315 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07438 313 316 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07437 8185 313 314 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07436 312 317 313 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07435 725 312 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07434 8185 312 725 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07433 4859 5022 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07432 4860 5023 5021 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07431 4858 5024 5017 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07430 8185 5015 4858 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07429 8185 5864 5024 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07428 5023 5024 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07427 8185 5027 5022 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07426 5021 5024 4859 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07425 5018 5021 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07424 8185 5018 4860 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07423 5017 5023 5018 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07422 5015 5017 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07421 8185 5017 5015 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07420 6630 6639 6631 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07419 6631 6629 6630 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07418 8185 6627 6631 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07417 7361 4955 4724 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07416 4724 4730 7361 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07415 8185 4731 4724 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07414 1280 2718 1281 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07413 1281 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07412 1279 4068 1280 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07411 1616 1394 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07410 1394 5648 1279 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07409 3501 3641 3502 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07408 3502 3642 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07407 3500 4299 3501 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07406 3660 3643 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07405 3643 4287 3500 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07404 447 5148 448 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07403 448 2203 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07402 446 1372 447 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07401 558 560 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07400 560 1157 446 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07399 252 254 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07398 251 253 250 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07397 247 255 248 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07396 8185 266 247 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07395 8185 1951 255 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07394 253 255 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07393 8185 256 254 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07392 250 255 252 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07391 249 250 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07390 8185 249 251 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07389 248 253 249 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07388 266 248 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07387 8185 248 266 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07386 8185 7314 7308 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07385 7160 7308 7307 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07384 8185 7513 7160 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07383 7484 7307 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07382 8185 7307 7484 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07381 7360 7791 7192 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07380 7192 7788 7360 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07379 8185 7824 7192 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07378 7358 7360 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07377 8185 2202 2412 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07376 2412 2198 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07375 8185 2199 2412 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07374 3009 2887 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07373 8185 2888 3009 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07372 3009 3606 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07371 8185 3603 3009 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07370 2140 2612 2046 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07369 2046 2141 2140 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07368 8185 2136 2046 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07367 2138 2140 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07366 7560 7562 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07365 7469 7470 7468 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07364 7466 7561 7557 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07363 8185 7558 7466 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07362 8185 7821 7561 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07361 7470 7561 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07360 8185 8139 7562 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07359 7468 7561 7560 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07358 7467 7468 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07357 8185 7467 7469 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07356 7557 7470 7467 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07355 7558 7557 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07354 8185 7557 7558 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07353 4812 6261 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07352 4885 8064 4812 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07351 6882 7110 6724 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07350 6724 7106 6882 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07349 8185 6880 6724 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07348 1216 4137 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07347 1490 1315 1216 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07346 7573 7576 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07345 7476 7477 7475 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07344 7473 7574 7570 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07343 8185 7572 7473 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07342 8185 8166 7574 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07341 7477 7574 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07340 8185 7575 7576 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07339 7475 7574 7573 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07338 7474 7475 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07337 8185 7474 7476 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07336 7570 7477 7474 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07335 7572 7570 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07334 8185 7570 7572 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07333 4323 4483 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07332 4322 4484 4482 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07331 4321 4485 4480 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07330 8185 7954 4321 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07329 8185 8063 4485 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07328 4484 4485 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07327 8185 7963 4483 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07326 4482 4485 4323 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07325 4481 4482 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07324 8185 4481 4322 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07323 4480 4484 4481 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07322 7954 4480 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07321 8185 4480 7954 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07320 8183 8179 8181 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07319 8181 8180 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07318 8182 8188 8183 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07317 7690 7884 7691 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07316 7691 7892 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07315 7890 7883 7690 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07314 835 2719 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07313 1154 2718 835 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07312 644 2719 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07311 1364 4067 644 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07310 8185 6363 3010 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07309 3010 3150 3151 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07308 3361 3151 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07307 4171 7029 4170 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07306 4170 5406 4171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07305 8185 6798 4170 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07304 8185 4492 3291 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07303 3291 3720 3290 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07302 3717 3290 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07301 6582 6585 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07300 6580 6584 6583 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07299 6578 6587 6577 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07298 8185 6576 6578 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07297 8185 7821 6587 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07296 6584 6587 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07295 8185 6581 6585 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07294 6583 6587 6582 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07293 6579 6583 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07292 8185 6579 6580 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07291 6577 6584 6579 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07290 6576 6577 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07289 8185 6577 6576 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07288 4367 7871 4571 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07287 8185 4571 4460 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07286 8185 7871 4464 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07285 4368 5030 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07284 4571 4464 4368 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07283 8185 4461 4367 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07282 4460 4571 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07281 6230 6383 6386 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07280 8185 6383 6384 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07279 6231 7622 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07278 6386 6384 6231 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07277 8185 6381 6230 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07276 2391 2408 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07275 2390 4433 2391 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07274 7651 7738 7650 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07273 7650 7729 7732 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07272 8185 7730 7651 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07271 7962 7732 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07270 8185 7343 7013 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07269 7013 7012 7014 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07268 7011 7014 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07267 8185 7759 7756 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07266 7659 7756 7755 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07265 8185 7753 7659 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07264 7754 7755 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07263 8185 7755 7754 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07262 8185 4032 3470 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07261 3470 3802 3607 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07260 3606 3607 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07259 2848 3327 2849 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07258 8185 2849 2847 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07257 8185 3327 2851 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07256 2850 3348 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07255 2849 2851 2850 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07254 8185 3315 2848 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_07253 2847 2849 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07252 7241 7310 7161 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07251 7161 7313 7241 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07250 8185 7311 7161 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07249 8185 7478 7220 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07248 7220 7405 7404 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07247 7304 7404 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07246 1966 1964 1967 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07245 1967 1965 1966 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07244 8185 4429 1967 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07243 8185 2256 2034 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07242 2034 2258 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07241 2039 2034 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07240 8185 2964 2967 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07239 2965 2967 2966 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07238 8185 2968 2965 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07237 3662 2966 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07236 8185 2966 3662 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07235 8185 3635 3637 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07234 3637 3636 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07233 4070 3637 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07232 2423 2430 2425 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07231 2425 2424 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07230 2422 2421 2423 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07229 2890 4203 2422 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07228 7499 7802 7498 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07227 7498 7747 7499 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07226 8185 7737 7498 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07225 7497 7499 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07224 4339 4574 4340 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07223 4340 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07222 4338 7051 4339 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07221 4424 5898 4338 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07220 5811 6658 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07219 5872 7151 5811 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07218 5810 6672 5872 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07217 8185 6668 5810 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07216 5810 6178 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_07215 3020 5942 3021 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07214 3021 5447 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07213 6363 7353 3020 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07212 8185 7137 5731 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07211 5731 5876 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07210 5730 5731 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07209 4927 1477 1478 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07208 1478 1476 4927 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07207 8185 3148 1478 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07206 1560 1559 1561 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07205 1561 1796 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07204 1557 1806 1560 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07203 1558 1556 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07202 1556 1891 1557 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07201 1883 5169 1884 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07200 1884 4517 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07199 1882 2227 1883 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07198 1985 1984 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07197 1984 4518 1882 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07196 2992 3106 3313 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07195 8185 3108 2992 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07194 2993 3109 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07193 3313 3107 2993 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07192 8185 3109 3106 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07191 3107 3108 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07190 6495 6278 6199 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07189 6199 6783 6495 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07188 8185 6279 6199 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07187 8185 3972 3887 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07186 3887 4648 3970 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07185 3969 3970 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07184 4521 4705 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07183 8185 8047 4521 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07182 4521 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07181 8185 8045 4521 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07180 4439 4521 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07179 8185 5132 5134 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07178 5134 5420 5135 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07177 5133 5135 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07176 8056 8064 8058 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07175 8185 8064 8062 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07174 8057 8059 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07173 8058 8062 8057 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07172 8185 8055 8056 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07171 8185 2492 768 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07170 768 1799 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07169 1800 768 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07168 8185 2962 2963 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07167 8185 3258 2963 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07166 2963 3865 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07165 2961 2963 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07164 8185 4068 2433 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07163 2433 6311 2432 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07162 2682 2432 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07161 8185 4945 4344 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07160 4344 4942 4519 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07159 4438 4519 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07158 8185 6302 6214 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07157 6214 6301 6303 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07156 6300 6303 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07155 8185 1996 1997 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07154 1997 1999 1998 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07153 2424 1998 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07152 8185 4167 2557 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07151 2557 4310 2691 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07150 3370 2691 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07149 4215 7354 4216 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07148 4216 4310 4217 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07147 8185 6293 4215 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07146 6089 4217 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07145 3875 3876 3874 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07144 3874 3872 3873 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07143 8185 4479 3875 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07142 3871 3873 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07141 4324 4487 4403 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07140 8185 4651 4324 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07139 4325 4489 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07138 4403 4488 4325 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07137 8185 4489 4487 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07136 4488 4651 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07135 3496 5447 3495 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07134 3495 7026 3634 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07133 8185 7353 3496 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07132 3842 3634 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_07131 8185 5940 388 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07130 388 2262 387 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07129 386 387 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07128 6800 6988 6696 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07127 6696 6835 6800 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07126 8185 7048 6696 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07125 6798 6800 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07124 1298 1293 1199 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07123 1199 1292 1298 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07122 8185 1954 1199 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07121 2498 2500 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07120 2497 2499 2496 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07119 2493 2501 2494 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07118 8185 2492 2493 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07117 8185 3834 2501 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07116 2499 2501 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07115 8185 3661 2500 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07114 2496 2501 2498 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07113 2495 2496 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07112 8185 2495 2497 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07111 2494 2499 2495 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07110 2492 2494 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07109 8185 2494 2492 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07108 6148 6149 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07107 6028 6030 6029 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07106 6026 6150 6144 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07105 8185 6145 6026 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07104 8185 7821 6150 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07103 6030 6150 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07102 8185 6617 6149 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07101 6029 6150 6148 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07100 6027 6029 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07099 8185 6027 6028 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07098 6144 6030 6027 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07097 6145 6144 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07096 8185 6144 6145 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07095 8185 5188 3616 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07094 7314 3616 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07093 8185 3616 7314 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07092 8185 3616 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07091 8144 3616 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07090 8185 5188 3808 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07089 8064 3808 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07088 8185 3808 8064 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07087 8185 3808 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07086 8144 3808 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07085 8185 5188 5172 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07084 7957 5172 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07083 8185 5172 7957 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07082 8185 5172 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07081 8144 5172 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07080 8185 5188 5173 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07079 7500 5173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07078 8185 5173 7500 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07077 8185 5173 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07076 8144 5173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07075 8185 4079 4080 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07074 5188 4080 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07073 8185 4080 5188 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07072 8185 4080 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07071 8144 4080 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07070 1684 4068 1685 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07069 1685 4575 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07068 1683 4167 1684 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07067 1825 1824 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07066 1824 7353 1683 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07065 2036 1827 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07064 8185 1825 2036 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07063 6667 6918 6664 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07062 6664 6663 6667 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07061 8185 7149 6664 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07060 1260 1372 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07059 8185 2698 1260 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07058 1260 4518 1821 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07057 1821 2926 1260 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07056 3459 3780 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07055 3581 5197 3459 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07054 331 330 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07053 328 332 329 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07052 326 333 325 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07051 8185 535 326 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07050 8185 3834 333 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07049 332 333 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07048 8185 549 330 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07047 329 333 331 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07046 327 329 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07045 8185 327 328 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07044 325 332 327 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07043 535 325 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07042 8185 325 535 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07041 7534 7779 7533 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07040 7533 7778 7534 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07039 8185 7585 7533 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07038 7783 7534 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07037 1602 4293 1603 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07036 1603 4310 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07035 1601 5483 1602 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07034 1898 1600 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_07033 1600 3857 1601 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07032 2864 2877 2865 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07031 2865 2866 2864 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07030 8185 2863 2865 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07029 3575 2864 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07028 4356 4546 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07027 4355 4547 4545 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07026 4354 4549 4542 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07025 8185 4543 4354 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07024 8185 5864 4549 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07023 4547 4549 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_07022 8185 5213 4546 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_07021 4545 4549 4356 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07020 4544 4545 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07019 8185 4544 4355 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07018 4542 4547 4544 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07017 4543 4542 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07016 8185 4542 4543 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07015 5145 7352 5146 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07014 5146 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07013 5144 5143 5145 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07012 6020 6359 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07011 6019 6363 6020 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07010 6613 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07009 7104 7095 6613 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07008 6608 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07007 6880 6870 6608 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_07006 3030 3787 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07005 8185 3787 3160 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_07004 8185 5453 3029 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07003 3161 3159 3030 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07002 3029 3160 3161 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07001 3158 3161 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_07000 8185 3161 3158 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06999 3159 5453 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06998 4277 5867 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06997 4276 4790 4277 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06996 8103 8106 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06995 8101 8105 8104 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06994 8098 8107 8099 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06993 8185 8097 8098 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06992 8185 8166 8107 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06991 8105 8107 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06990 8185 8102 8106 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06989 8104 8107 8103 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06988 8100 8104 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06987 8185 8100 8101 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06986 8099 8105 8100 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06985 8097 8099 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06984 8185 8099 8097 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06983 5311 5629 5312 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06982 5312 5628 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06981 6480 5434 5311 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06980 6033 7872 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06979 6400 6652 6033 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06978 742 903 741 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06977 8185 741 740 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06976 8185 903 744 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06975 743 4176 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06974 741 744 743 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06973 8185 739 742 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06972 740 741 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06971 4177 4178 4179 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06970 8185 4179 4176 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06969 8185 4178 4181 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06968 4180 4925 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06967 4179 4181 4180 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06966 8185 8139 4177 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06965 4176 4179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06964 4638 7887 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06963 4786 7130 4638 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06962 3846 3857 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06961 3847 3844 3846 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06960 3845 4575 3847 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06959 8185 7788 3845 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06958 3845 3842 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06957 3912 4517 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06956 4010 4518 3912 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06955 8185 4009 4010 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06954 4192 4010 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06953 1926 2152 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06952 1927 2608 1926 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06951 8185 2616 1927 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06950 1925 1927 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06949 8185 4512 3901 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06948 3901 4511 3992 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06947 3991 3992 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06946 3134 1760 1653 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06945 1653 1761 3134 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06944 8185 1962 1653 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06943 3005 4172 3006 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06942 3006 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06941 3146 8122 3005 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06940 2862 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06939 2875 3139 2862 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06938 2861 3130 2875 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06937 8185 3737 2861 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06936 2861 2860 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06935 6481 6524 5745 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06934 5745 6294 6481 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06933 8185 5886 5745 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06932 5588 5414 5296 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06931 5296 5616 5588 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06930 8185 7957 5296 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06929 7623 7883 7625 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06928 7624 7627 7623 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06927 7625 7884 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06926 7622 7623 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06925 8185 7876 7624 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06924 7624 7877 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06923 5798 7126 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06922 5858 6154 5798 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06921 1225 1332 1334 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06920 8185 1334 1330 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06919 8185 1332 1336 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06918 1226 4012 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06917 1334 1336 1226 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06916 8185 1335 1225 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06915 1330 1334 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06914 1075 1332 1077 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06913 8185 1077 1074 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06912 8185 1332 1078 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06911 1076 4160 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06910 1077 1078 1076 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06909 8185 1317 1075 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06908 1074 1077 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06907 3022 7026 3023 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06906 3023 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06905 4548 6796 3022 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06904 3019 6543 3018 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06903 3018 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06902 5434 6544 3019 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06901 1569 7026 1568 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06900 1568 6543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06899 1887 4293 1569 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06898 6751 7643 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06897 6920 7869 6751 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06896 3950 4068 3949 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06895 3949 4295 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06894 3948 7026 3950 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06893 4298 4067 3948 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06892 4381 4790 4380 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06891 4380 6421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06890 4379 7887 4381 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06889 4473 5740 4379 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06888 4390 4517 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06887 6286 4518 4390 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06886 8185 7957 7961 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06885 7958 7961 7959 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06884 8185 8008 7958 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06883 7956 7959 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06882 8185 7959 7956 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06881 3821 5447 3820 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06880 3820 4574 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06879 3818 6293 3821 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06878 3819 4260 3818 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06877 8185 2159 2058 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06876 2058 5401 2160 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06875 2619 2160 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06874 8185 2866 2542 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06873 2542 2877 2658 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06872 2659 2658 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06871 7230 7338 7231 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06870 7231 7340 7337 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06869 8185 7339 7230 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06868 7332 7337 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06867 7224 7725 7223 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06866 7223 7749 7315 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06865 8185 7724 7224 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06864 7313 7315 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06863 1221 1332 1323 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06862 8185 1323 1506 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06861 8185 1332 1324 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06860 1222 4176 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06859 1323 1324 1222 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06858 8185 1499 1221 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06857 1506 1323 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06856 717 1332 918 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06855 8185 918 915 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06854 8185 1332 919 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06853 719 3999 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06852 918 919 719 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06851 8185 1088 717 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06850 915 918 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06849 1092 1332 1094 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06848 8185 1094 1091 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06847 8185 1332 1096 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06846 1093 2402 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06845 1094 1096 1093 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06844 8185 1758 1092 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06843 1091 1094 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06842 695 939 897 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06841 8185 897 1069 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06840 8185 939 898 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06839 696 3537 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06838 897 898 696 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06837 8185 1063 695 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06836 1069 897 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06835 275 939 274 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06834 8185 274 272 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06833 8185 939 277 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06832 276 3532 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06831 274 277 276 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06830 8185 273 275 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06829 272 274 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06828 3016 4574 3017 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06827 3017 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06826 5169 6293 3016 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06825 8185 1593 1594 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06824 1594 1597 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06823 1892 1594 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06822 8185 3556 2820 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06821 2817 2813 2814 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06820 2821 3757 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_06819 2814 2815 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06818 8185 3556 2815 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_06817 3095 2817 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_06816 2820 2816 2818 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06815 2818 3757 2817 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06814 2817 2821 2819 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06813 2819 3303 2820 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06812 8185 3556 2522 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06811 2626 2619 2519 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06810 2623 3757 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_06809 2519 2620 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06808 8185 3556 2620 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_06807 3098 2626 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_06806 2522 2621 2520 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06805 2520 3757 2626 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06804 2626 2623 2521 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06803 2521 3307 2522 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_06802 5647 5908 5646 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06801 5646 6359 5645 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06800 8185 6363 5647 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06799 5644 5645 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06798 404 939 502 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06797 8185 502 691 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06796 8185 939 456 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06795 405 3978 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06794 502 456 405 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06793 8185 685 404 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06792 691 502 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06791 745 939 937 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06790 8185 937 935 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06789 8185 939 940 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06788 746 4012 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06787 937 940 746 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06786 8185 1113 745 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06785 935 937 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06784 1562 4572 1563 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06783 1563 4573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06782 1796 4574 1562 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06781 6184 7893 6183 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06780 6183 8187 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06779 6182 6893 6184 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06778 6189 7883 6182 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06777 4809 6636 4808 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06776 4808 5875 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06775 4807 6396 4809 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06774 5041 6921 4807 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06773 5274 6172 5275 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06772 5275 6652 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06771 5272 6421 5274 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06770 5273 6921 5272 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06769 4393 4529 4392 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06768 4392 4707 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06767 4391 4548 4393 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06766 7761 4524 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06765 4524 4527 4391 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06764 8185 4766 4768 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06763 4768 5501 4767 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06762 4765 4767 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06761 8185 7880 4853 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06760 4853 5701 5001 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06759 5002 5001 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06758 8185 8064 1124 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06757 1124 1132 1125 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06756 1123 1125 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06755 7800 7802 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06754 8185 8047 7800 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06753 7800 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06752 8185 8045 7800 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06751 7801 7800 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06750 3454 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06749 3570 3571 3454 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06748 3453 3569 3570 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06747 8185 3737 3453 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06746 3453 3567 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06745 6208 6775 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06744 6290 6480 6208 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06743 8185 6295 6290 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06742 6500 6290 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06741 8185 4556 4360 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06740 4360 6383 4555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06739 5212 4555 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06738 8185 370 183 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06737 4310 183 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06736 8185 183 4310 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06735 8185 183 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06734 8144 183 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06733 8185 370 371 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06732 1565 371 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06731 8185 371 1565 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06730 8185 371 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06729 8144 371 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06728 8185 185 182 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06727 370 182 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06726 8185 182 370 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06725 8185 182 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06724 8144 182 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06723 8185 1968 1763 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06722 8045 1763 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06721 8185 1763 8045 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06720 8185 1763 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06719 8144 1763 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06718 8185 1968 1969 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06717 4429 1969 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06716 8185 1969 4429 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06715 8185 1969 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06714 8144 1969 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06713 8185 1776 1764 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06712 1968 1764 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06711 8185 1764 1968 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06710 8185 1764 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06709 8144 1764 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06708 8185 5654 2910 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06707 2910 4167 2911 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06706 3371 2911 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06705 1326 1327 1223 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06704 1223 1325 1326 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06703 8185 1962 1223 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06702 3997 1326 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06701 6194 6267 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06700 6268 6480 6194 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06699 8185 6266 6268 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06698 6472 6268 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06697 4237 4236 4238 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06696 4238 6867 4237 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06695 8185 7867 4238 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06694 4738 4237 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06693 2426 4067 2428 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06692 2427 6796 2426 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06691 2428 2896 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06690 2677 2426 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06689 8185 2898 2427 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06688 2427 2894 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06687 7585 7280 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06686 7528 7073 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06685 8185 8184 6646 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06684 6646 7884 6649 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06683 6663 6649 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06682 2584 4575 2585 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06681 2585 4310 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06680 2583 4302 2584 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06679 2950 2725 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06678 2725 5483 2583 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06677 1247 1996 1246 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06676 1246 4540 1363 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06675 8185 1986 1247 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06674 1362 1363 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06673 356 1150 355 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06672 355 359 357 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06671 8185 4251 356 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06670 354 357 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06669 1911 6469 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06668 1912 7728 1911 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06667 8185 1909 1912 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06666 1910 1912 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06665 2524 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06664 3109 2836 2524 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06663 2523 3112 3109 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06662 8185 3737 2523 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06661 2523 3108 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06660 283 284 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06659 281 285 282 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06658 279 286 278 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06657 8185 512 279 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06656 8185 1951 286 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06655 285 286 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06654 8185 287 284 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06653 282 286 283 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06652 280 282 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06651 8185 280 281 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06650 278 285 280 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06649 512 278 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06648 8185 278 512 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06647 3940 4059 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06646 3941 4060 4058 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06645 3939 4062 4054 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06644 8185 4461 3939 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06643 8185 5864 4062 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06642 4060 4062 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06641 8185 4460 4059 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06640 4058 4062 3940 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06639 4055 4058 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06638 8185 4055 3941 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06637 4054 4060 4055 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06636 4461 4054 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06635 8185 4054 4461 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06634 4330 4500 4414 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06633 8185 5109 4330 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06632 4331 4672 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06631 4414 4501 4331 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06630 8185 4672 4500 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06629 4501 5109 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06628 844 6609 843 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06627 843 4068 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06626 842 4306 844 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06625 1168 960 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06624 960 3857 842 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06623 7349 7061 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06622 3945 5483 3946 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06621 3946 5447 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06620 3944 7051 3945 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06619 4790 4064 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06618 4064 4075 3944 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06617 3770 4939 3769 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06616 3769 5406 3770 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06615 8185 6553 3769 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06614 3768 3770 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06613 2598 2596 2506 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06612 2506 3287 2598 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06611 8185 2594 2506 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06610 2595 2598 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06609 398 492 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06608 397 493 491 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06607 396 494 486 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06606 8185 497 396 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06605 8185 1951 494 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06604 493 494 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06603 8185 496 492 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06602 491 494 398 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06601 489 491 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06600 8185 489 397 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06599 486 493 489 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06598 497 486 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06597 8185 486 497 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06596 7678 7842 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06595 7679 7843 7841 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06594 7677 7844 7837 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06593 8185 7835 7677 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06592 8185 8166 7844 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06591 7843 7844 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06590 8185 7863 7842 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06589 7841 7844 7678 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06588 7838 7841 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06587 8185 7838 7679 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06586 7837 7843 7838 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06585 7835 7837 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06584 8185 7837 7835 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06583 1880 4184 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06582 1978 1966 1880 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06581 4291 4295 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06580 4292 4997 4291 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06579 4290 4790 4292 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06578 8185 5732 4290 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06577 4290 6912 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_06576 7682 7853 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06575 7681 7854 7849 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06574 7680 7855 7846 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06573 8185 7845 7680 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06572 8185 8166 7855 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06571 7854 7855 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06570 8185 7851 7853 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06569 7849 7855 7682 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06568 7848 7849 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06567 8185 7848 7681 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06566 7846 7854 7848 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06565 7845 7846 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06564 8185 7846 7845 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06563 2503 6472 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06562 6083 6473 2503 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06561 2547 2677 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06560 2678 6076 2547 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06559 7548 2492 363 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06558 8185 1799 364 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06557 363 364 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06556 1237 1558 1238 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06555 1238 1357 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06554 1962 1355 1237 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06553 3317 3748 3319 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06552 8185 3319 3316 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06551 8185 3748 3321 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06550 3318 3348 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06549 3319 3321 3318 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06548 8185 3315 3317 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06547 3316 3319 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06546 391 474 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06545 392 475 472 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06544 390 476 469 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06543 8185 3077 390 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06542 8185 3708 476 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06541 475 476 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06540 8185 1910 474 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06539 472 476 391 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06538 470 472 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06537 8185 470 392 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06536 469 475 470 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06535 3077 469 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06534 8185 469 3077 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06533 8185 7343 7039 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06532 7039 7048 7040 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06531 7038 7040 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06530 8001 8094 8003 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06529 8185 8003 7999 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06528 8185 8094 8005 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06527 8002 8015 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06526 8003 8005 8002 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06525 8185 8000 8001 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06524 7999 8003 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06523 8022 8094 8023 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06522 8185 8023 8020 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06521 8185 8094 8027 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06520 8024 8038 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06519 8023 8027 8024 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06518 8185 8021 8022 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06517 8020 8023 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06516 8041 8094 8042 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06515 8185 8042 8039 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06514 8185 8094 8044 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06513 8043 8066 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06512 8042 8044 8043 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06511 8185 8040 8041 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06510 8039 8042 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06509 8088 8094 8087 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06508 8185 8087 8085 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06507 8185 8094 8091 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06506 8090 8089 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06505 8087 8091 8090 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06504 8185 8086 8088 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06503 8085 8087 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06502 8072 8094 8074 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06501 8185 8074 8070 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06500 8185 8094 8075 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06499 8073 8109 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06498 8074 8075 8073 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06497 8185 8071 8072 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06496 8070 8074 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06495 7567 8094 7569 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06494 8185 7569 7829 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06493 8185 8094 7571 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06492 7568 8136 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06491 7569 7571 7568 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06490 8185 7824 7567 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06489 7829 7569 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06488 631 3711 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06487 3063 1047 631 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06486 4701 4714 4621 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06485 8185 7314 4622 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06484 4621 4622 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06483 562 1799 450 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06482 8185 2492 563 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06481 450 563 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06480 8185 2477 2026 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06479 2023 2026 2024 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06478 8185 2022 2023 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06477 2238 2024 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06476 8185 2024 2238 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06475 2080 2206 2079 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06474 2079 2207 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06473 2888 2205 2080 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06472 8185 3553 2048 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06471 2048 2803 2142 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06470 2141 2142 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06469 4333 5648 4334 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06468 4334 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06467 4332 7051 4333 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06466 4512 6489 4332 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06465 2320 3752 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06464 2319 2318 2320 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06463 6686 6784 6685 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06462 6685 6786 6787 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06461 8185 6785 6686 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06460 6783 6787 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06459 8092 8094 8093 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06458 8185 8093 8102 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06457 8185 8094 8096 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06456 8095 8156 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06455 8093 8096 8095 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06454 8185 8097 8092 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06453 8102 8093 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06452 5702 7872 5703 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06451 5703 8179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06450 5700 7633 5702 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06449 5701 7130 5700 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06448 821 1154 822 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06447 822 4228 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06446 820 5147 821 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06445 1358 954 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06444 954 1543 820 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06443 3927 4572 3929 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06442 3929 7354 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06441 3928 5447 3927 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06440 4234 4031 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06439 4031 6143 3928 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06438 8185 3997 3998 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06437 3905 3998 3996 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06436 8185 4690 3905 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06435 3995 3996 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06434 8185 3996 3995 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06433 6475 6478 6479 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06432 6479 6477 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06431 6476 6472 6475 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06430 7724 6474 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06429 6474 6473 6476 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06428 6055 7029 5751 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06427 5751 6294 6055 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06426 8185 5897 5751 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06425 8185 7056 5116 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06424 5116 5114 5115 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06423 5113 5115 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06422 8185 2262 186 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06421 56 186 184 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06420 8185 5940 56 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06419 185 184 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06418 8185 184 185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06417 7696 7893 7697 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06416 7697 7892 7894 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06415 8185 7891 7696 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06414 8180 7894 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06413 8185 1758 1652 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06412 1652 5641 1759 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06411 2178 1759 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06410 8185 1499 1220 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06409 1220 5641 1320 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06408 1964 1320 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06407 4151 4153 4152 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06406 8185 4149 4151 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06405 4154 4498 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06404 4152 4150 4154 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06403 8185 4498 4153 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06402 4150 4149 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06401 8185 4129 4131 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06400 4131 4133 4132 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06399 4130 4132 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06398 8185 4734 3402 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06397 3402 4075 3403 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06396 3399 3403 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06395 2913 4306 2558 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06394 2558 4302 2913 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06393 8185 3371 2558 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06392 5402 7020 5294 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06391 5294 5406 5402 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06390 8185 6788 5294 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06389 5401 5402 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06388 1648 1749 4489 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06387 8185 6793 1648 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06386 1649 4402 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06385 4489 1750 1649 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06384 8185 4402 1749 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06383 1750 6793 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06382 6746 7881 6747 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06381 6747 7403 6913 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06380 8185 7891 6746 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06379 6918 6913 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06378 3862 4476 3861 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06377 3861 3863 3864 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06376 8185 4299 3862 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06375 3860 3864 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06374 3422 3425 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06373 3272 3424 3271 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06372 3269 3426 3421 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06371 8185 5940 3269 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06370 8185 3834 3426 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06369 3424 3426 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06368 8185 3423 3425 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06367 3271 3426 3422 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06366 3270 3271 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06365 8185 3270 3272 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06364 3421 3424 3270 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06363 5940 3421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06362 8185 3421 5940 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06361 8185 7957 5548 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06360 5547 5548 5549 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06359 8185 7752 5547 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06358 7481 5549 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06357 8185 5549 7481 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06356 4758 6412 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06355 4757 5002 4758 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06354 8185 4756 4757 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06353 7355 7791 7191 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06352 7191 7788 7355 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06351 8185 8086 7191 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06350 7257 7355 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06349 2108 2247 2109 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06348 2109 2246 2248 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06347 8185 3172 2108 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06346 2958 2248 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06345 1177 6609 1178 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06344 1178 4068 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06343 1176 6796 1177 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06342 1173 1175 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06341 1175 3857 1176 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06340 4785 7130 4784 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06339 4784 7887 4783 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06338 8185 7149 4785 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06337 4782 4783 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06336 338 344 340 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06335 340 352 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06334 339 551 338 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06333 5641 337 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06332 337 349 339 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06331 8185 3340 2867 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06330 2867 3009 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06329 2866 2867 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06328 5218 5222 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06327 5220 5221 5219 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06326 5215 5224 5216 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06325 8185 5485 5215 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06324 8185 5864 5224 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06323 5221 5224 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06322 8185 5490 5222 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06321 5219 5224 5218 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06320 5217 5219 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06319 8185 5217 5220 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06318 5216 5221 5217 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06317 5485 5216 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06316 8185 5216 5485 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06315 1689 5447 1690 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06314 1690 4067 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06313 1688 5942 1689 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06312 1904 1829 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06311 1829 4075 1688 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06310 23 120 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06309 22 121 119 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06308 21 122 115 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06307 8185 514 21 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06306 8185 1951 122 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06305 121 122 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06304 8185 292 120 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06303 119 122 23 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06302 116 119 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06301 8185 116 22 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06300 115 121 116 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06299 514 115 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06298 8185 115 514 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06297 5331 5464 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06296 5330 5465 5463 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06295 5329 5466 5459 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06294 8185 5670 5329 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06293 8185 7821 5466 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06292 5465 5466 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06291 8185 5671 5464 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06290 5463 5466 5331 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06289 5460 5463 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06288 8185 5460 5330 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06287 5459 5465 5460 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06286 5670 5459 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06285 8185 5459 5670 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06284 3706 3707 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06283 3704 3710 3705 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06282 3702 3709 3701 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06281 8185 3956 3702 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06280 8185 3708 3709 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06279 3710 3709 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06278 8185 3955 3707 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06277 3705 3709 3706 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06276 3703 3705 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06275 8185 3703 3704 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06274 3701 3710 3703 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06273 3956 3701 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06272 8185 3701 3956 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06271 4629 4737 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06270 8140 4739 4629 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06269 6239 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06268 6399 6398 6239 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06267 5711 6654 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06266 5710 6652 5711 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06265 3506 3877 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06264 3667 4318 3506 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06263 7655 7741 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06262 7740 7743 7655 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06261 8185 7744 7740 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06260 7985 7740 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06259 4033 4770 3930 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06258 8185 6143 4034 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06257 3930 4034 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06256 2067 3348 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06255 3229 3315 2067 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06254 6545 6543 6546 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06253 6546 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06252 6542 6544 6545 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06251 7338 6541 6542 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06250 1135 5654 1136 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06249 1136 5648 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06248 1356 1353 1135 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06247 6730 7297 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06246 6899 6897 6730 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06245 5799 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06244 5862 6141 5799 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06243 4637 6383 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06242 5223 5003 4637 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06241 415 903 527 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06240 8185 527 528 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06239 8185 903 459 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06238 416 3999 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06237 527 459 416 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06236 8185 517 415 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06235 528 527 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06234 2562 6543 2561 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06233 2561 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06232 6359 4293 2562 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06231 7479 8186 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06230 7478 8184 7479 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06229 4398 6191 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06228 4479 4790 4398 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06227 8185 2032 1899 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06226 1899 1821 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06225 8185 2249 1899 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06224 5149 5147 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06223 6285 5148 5149 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06222 1206 5395 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06221 2144 1301 1206 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06220 2396 2400 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06219 2395 2399 2397 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06218 2392 2401 2393 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06217 8185 6080 2392 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06216 8185 3708 2401 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06215 2399 2401 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_06214 8185 2398 2400 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_06213 2397 2401 2396 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06212 2394 2397 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06211 8185 2394 2395 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06210 2393 2399 2394 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06209 6080 2393 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06208 8185 2393 6080 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06207 7164 7749 7165 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06206 7165 7518 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06205 7163 7725 7164 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06204 7490 7724 7163 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06203 7320 7766 7169 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06202 7169 7747 7320 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06201 8185 7748 7169 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06200 7316 7320 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06199 3906 4178 4002 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06198 8185 4002 3999 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06197 8185 4178 4004 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06196 3907 4698 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06195 4002 4004 3907 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06194 8185 7863 3906 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06193 3999 4002 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06192 30 903 144 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06191 8185 144 141 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06190 8185 903 145 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06189 31 2402 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06188 144 145 31 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06187 8185 530 30 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06186 141 144 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06185 4504 4507 4389 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06184 4388 7550 4504 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06183 4389 4701 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06182 4418 4504 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06181 8185 7548 4388 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06180 4388 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06179 3475 4051 3476 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06178 3476 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06177 4527 4067 3475 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06176 7554 7558 7462 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06175 8185 7957 7463 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06174 7462 7463 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06173 3490 5648 3489 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06172 3489 6543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06171 3488 6544 3490 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06170 3625 3857 3488 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06169 3493 6797 3494 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06168 3494 4295 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06167 3492 7026 3493 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06166 3628 6544 3492 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06165 3866 4474 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06164 3865 4311 3866 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06163 3259 4292 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06162 3258 4468 3259 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06161 8185 5453 2548 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06160 2548 2679 2680 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06159 2887 2680 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06158 8185 4166 2837 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06157 2837 3759 2839 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06156 2836 2839 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06155 8185 3134 3001 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06154 3001 4947 3136 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06153 3135 3136 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06152 8185 3229 2534 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06151 2534 2868 2647 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06150 2853 2647 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06149 6032 6906 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06148 6157 6905 6032 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06147 711 939 713 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06146 8185 713 710 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06145 8185 939 714 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06144 712 4160 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06143 713 714 712 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06142 8185 709 711 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06141 710 713 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06140 426 939 548 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06139 8185 548 549 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06138 8185 939 462 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06137 427 4176 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06136 548 462 427 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06135 8185 535 426 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06134 549 548 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06133 293 939 294 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06132 8185 294 292 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06131 8185 939 296 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06130 295 3999 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06129 294 296 295 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06128 8185 514 293 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06127 292 294 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06126 321 939 322 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06125 8185 322 320 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06124 8185 939 324 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06123 323 2402 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06122 322 324 323 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06121 8185 532 321 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06120 320 322 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06119 2404 5148 2403 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06118 8185 2403 2402 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06117 8185 5148 2406 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06116 2405 8122 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06115 2403 2406 2405 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06114 8185 6076 2404 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06113 2402 2403 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06112 1146 5148 1147 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06111 1147 4540 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06110 1144 1996 1146 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06109 1145 1372 1144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06108 5139 7787 5128 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06107 5128 5907 5139 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06106 8185 6549 5128 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06105 2107 2935 2106 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06104 2106 2240 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06103 2941 2462 2107 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06102 1741 1761 1495 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06101 1495 1760 1741 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06100 8185 3148 1495 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06099 6210 7356 6211 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06098 6211 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06097 6209 6293 6210 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06096 7002 6292 6209 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06095 3895 4172 3894 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06094 3894 4173 3988 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06093 8185 7349 3895 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06092 3987 3988 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06091 5305 5424 5304 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06090 5304 5428 5425 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06089 8185 5619 5305 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06088 5911 5425 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06087 4395 4548 4394 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06086 4394 4529 4528 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06085 8185 4527 4395 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06084 6294 4528 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_06083 673 903 672 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06082 8185 672 671 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06081 8185 903 675 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06080 674 3537 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06079 672 675 674 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06078 8185 677 673 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06077 671 672 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06076 3302 4178 3540 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06075 8185 3540 3537 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06074 8185 4178 3541 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06073 3304 4662 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06072 3540 3541 3304 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06071 8185 7549 3302 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_06070 3537 3540 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06069 6985 6992 6984 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06068 8185 7957 6986 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06067 6984 6986 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06066 4220 5654 4221 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06065 4221 4574 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06064 4219 6293 4220 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06063 4503 4218 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06062 4218 5938 4219 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06061 7878 7876 7686 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06060 7686 7877 7878 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06059 8185 7889 7686 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06058 3886 5453 3885 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06057 3885 6520 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06056 3884 5938 3886 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06055 3968 5606 3884 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06054 8185 4439 4201 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06053 4201 5150 4200 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06052 4198 4200 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06051 3004 3146 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06050 3144 4007 3004 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06049 8185 4510 3144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06048 3145 3144 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06047 5587 5898 5295 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06046 8185 8064 5404 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06045 5295 5404 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06044 7128 7884 7127 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06043 7129 7877 7128 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06042 7127 7869 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06041 7126 7128 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06040 8185 7885 7129 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06039 7129 7296 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_06038 8185 6793 5278 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06037 5278 5383 5378 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06036 5377 5378 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06035 3163 3171 3031 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06034 3031 3170 3163 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06033 8185 4742 3031 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06032 3250 3163 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06031 3632 4071 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06030 8185 3635 3632 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06029 3632 3629 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06028 8185 3636 3632 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06027 3651 3632 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06026 8185 1088 1090 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06025 1090 5641 1089 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06024 1760 1089 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06023 8185 1048 1049 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06022 1049 5641 1050 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06021 1476 1050 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06020 5666 7352 5668 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06019 8185 7352 5669 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06018 5667 6359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06017 5668 5669 5667 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06016 8185 6358 5666 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06015 7124 7888 7125 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06014 7125 7619 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06013 7122 8187 7124 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06012 7121 7123 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_06011 7123 8184 7122 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_06010 8185 4540 2096 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_06009 2096 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_06008 2234 2226 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06007 2096 7343 2226 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_06006 2226 2926 2096 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_06005 6595 6601 6598 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06004 8185 6594 6595 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06003 6599 6597 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06002 6598 6596 6599 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_06001 8185 6597 6601 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_06000 6596 6594 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05999 8185 4518 2880 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05998 2880 4517 2881 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05997 4203 2881 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05996 2181 2178 2068 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05995 2068 2179 2181 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05994 8185 4429 2068 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05993 554 1798 431 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05992 431 7548 554 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05991 8185 6363 431 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05990 557 554 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05989 2886 7779 2885 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05988 2885 7778 2886 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05987 8185 8122 2885 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05986 7539 8051 7538 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05985 7540 7550 7539 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05984 7538 8061 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05983 7536 7539 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05982 8185 7548 7540 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05981 7540 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05980 1564 6609 1566 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05979 1566 1565 1567 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05978 8185 4306 1564 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05977 4178 1567 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05976 1641 2346 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05975 1727 2610 1641 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05974 8185 2616 1727 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05973 4189 4939 4190 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05972 4190 5406 4189 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05971 8185 6553 4190 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05970 5569 5567 5568 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05969 5568 5633 5569 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05968 8185 6763 5568 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05967 5566 5569 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05966 1907 5648 1908 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05965 1908 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05964 1906 4067 1907 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05963 2043 2042 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05962 2042 5447 1906 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05961 8139 7612 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05960 7777 6988 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05959 4868 6396 4869 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05958 4869 5875 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05957 4867 6172 4868 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05956 5032 5033 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05955 5033 6921 4867 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05954 5733 6921 5735 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05953 5735 6914 5734 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05952 8185 7130 5733 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05951 5732 5734 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05950 270 1115 271 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05949 271 1114 269 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05948 269 273 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05947 267 266 271 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05946 8185 1110 267 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05945 8185 268 270 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05944 1744 271 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05943 2083 2430 2084 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05942 2084 2424 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05941 2082 2421 2083 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05940 2407 2209 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05939 2209 4203 2082 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05938 4147 4152 4148 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05937 4148 4416 4147 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05936 8185 4156 4148 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05935 4492 4147 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05934 26 129 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05933 25 130 126 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05932 24 131 123 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05931 8185 529 24 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05930 8185 1772 131 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05929 130 131 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05928 8185 306 129 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05927 126 131 26 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05926 125 126 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05925 8185 125 25 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05924 123 130 125 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05923 529 123 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05922 8185 123 529 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05921 4363 4561 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05920 4362 4562 4560 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05919 4361 4563 4557 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05918 8185 4558 4361 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05917 8185 5864 4563 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05916 4562 4563 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05915 8185 4765 4561 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05914 4560 4563 4363 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05913 4559 4560 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05912 8185 4559 4362 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05911 4557 4562 4559 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05910 4558 4557 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05909 8185 4557 4558 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05908 7535 7779 7537 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05907 7537 7778 7535 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05906 8185 7549 7537 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05905 7768 7535 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05904 1525 4025 1524 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05903 1524 1778 1525 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05902 8185 4198 1524 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05901 2540 2875 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05900 2863 2873 2540 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05899 735 737 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05898 639 736 732 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05897 638 738 730 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05896 8185 1111 638 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05895 8185 1772 738 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05894 736 738 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05893 8185 920 737 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05892 732 738 735 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05891 733 732 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05890 8185 733 639 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05889 730 736 733 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05888 1111 730 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05887 8185 730 1111 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05886 7362 7779 7193 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05885 7193 7778 7362 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05884 8185 8139 7193 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05883 7357 7362 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05882 1498 5136 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05881 1530 1497 1498 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05880 3239 4573 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05879 7559 7026 3239 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05878 7406 4024 3920 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05877 3920 4025 7406 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05876 8185 4207 3920 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05875 6555 8058 6556 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05874 6556 6835 6555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05873 8185 6554 6556 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05872 6553 6555 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05871 2535 2868 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05870 2652 3229 2535 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05869 7670 7811 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05868 7669 7812 7810 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05867 7668 7813 7806 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05866 8185 8059 7668 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05865 8185 8063 7813 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05864 7812 7813 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05863 8185 8122 7811 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05862 7810 7813 7670 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05861 7807 7810 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05860 8185 7807 7669 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05859 7806 7812 7807 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05858 8059 7806 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05857 8185 7806 8059 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05856 5 70 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05855 4 71 69 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05854 3 72 65 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05853 8185 6484 3 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05852 8185 1951 72 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05851 71 72 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05850 8185 3511 70 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05849 69 72 5 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05848 67 69 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05847 8185 67 4 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05846 65 71 67 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05845 6484 65 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05844 8185 65 6484 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05843 3349 8064 3588 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05842 8185 3588 3596 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05841 8185 8064 3591 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05840 3352 3787 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05839 3588 3591 3352 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05838 8185 4712 3349 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05837 3596 3588 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05836 7135 7158 7134 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05835 7134 7877 7135 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05834 8185 7885 7134 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05833 6421 8187 6258 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05832 6258 7893 6421 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05831 8185 7869 6258 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05830 3858 4798 3859 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05829 3859 3856 3858 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05828 8185 3857 3859 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05827 418 1115 534 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05826 534 1114 419 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05825 419 532 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05824 417 529 534 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05823 8185 1110 417 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05822 8185 530 418 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05821 2179 534 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05820 7178 7352 7179 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05819 7179 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05818 7327 8040 7178 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05817 1989 4572 1990 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05816 1990 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05815 2206 2968 1989 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05814 7205 7383 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05813 7204 7385 7381 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05812 7203 7382 7378 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05811 8185 7379 7203 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05810 8185 8166 7382 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05809 7385 7382 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05808 8185 7384 7383 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05807 7381 7382 7205 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05806 7380 7381 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05805 8185 7380 7204 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05804 7378 7385 7380 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05803 7379 7378 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05802 8185 7378 7379 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05801 6675 6759 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05800 6676 6760 6758 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05799 6674 6761 6754 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05798 8185 7513 6674 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05797 8185 8063 6761 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05796 6760 6761 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05795 8185 7485 6759 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05794 6758 6761 6675 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05793 6755 6758 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05792 8185 6755 6676 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05791 6754 6760 6755 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05790 7513 6754 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05789 8185 6754 7513 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05788 1976 8094 2194 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05787 8185 2194 2398 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05786 8185 8094 2196 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05785 1977 2390 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05784 2194 2196 1977 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05783 8185 6080 1976 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05782 2398 2194 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05781 2983 8094 3092 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05780 8185 3092 3282 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05779 8185 8094 3065 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05778 2984 3063 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05777 3092 3065 2984 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05776 8185 5563 2983 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05775 3282 3092 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05774 3299 8094 3298 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05773 8185 3298 3519 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05772 8185 8094 3301 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05771 3297 3300 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05770 3298 3301 3297 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05769 8185 5387 3299 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05768 3519 3298 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05767 1212 8094 1309 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05766 8185 1309 1307 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05765 8185 8094 1311 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05764 1213 1474 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05763 1309 1311 1213 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05762 8185 5394 1212 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05761 1307 1309 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05760 1520 8094 1521 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05759 8185 1521 1519 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05758 8185 8094 1523 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05757 1522 1525 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05756 1521 1523 1522 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05755 8185 5419 1520 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05754 1519 1521 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05753 1489 8094 1492 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05752 8185 1492 1488 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05751 8185 8094 1493 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05750 1491 1490 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05749 1492 1493 1491 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05748 8185 5571 1489 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05747 1488 1492 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05746 5107 5938 5106 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05745 5106 5108 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05744 5114 5606 5107 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05743 1051 2805 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05742 3300 1052 1051 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05741 449 4310 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05740 764 5483 449 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05739 8185 3315 1946 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05738 1946 3348 1945 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05737 2616 1945 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05736 8185 3542 1921 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05735 1921 2796 1920 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05734 2135 1920 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05733 8185 4543 3775 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05732 3775 3780 3777 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05731 3774 3777 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05730 3440 3990 3439 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05729 3439 3989 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05728 3438 3586 3440 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05727 3543 3581 3438 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05726 2661 2877 2541 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05725 2541 2866 2661 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05724 8185 7314 2541 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05723 1975 8094 1979 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05722 8185 1979 1974 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05721 8185 8094 1980 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05720 1981 1978 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05719 1979 1980 1981 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05718 8185 5435 1975 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05717 1974 1979 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05716 1527 8094 1529 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05715 8185 1529 1526 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05714 8185 8094 1531 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05713 1528 1530 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05712 1529 1531 1528 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05711 8185 5443 1527 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05710 1526 1529 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05709 1971 8094 1970 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05708 8185 1970 2189 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05707 8185 8094 1972 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05706 1973 2182 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05705 1970 1972 1973 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05704 8185 5143 1971 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05703 2189 1970 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05702 3925 4572 3926 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05701 3926 7354 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05700 3924 5447 3925 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05699 4725 6143 3924 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05698 4129 7787 3280 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05697 3280 5907 4129 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05696 8185 6292 3280 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05695 1497 1760 1496 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05694 1496 1761 1497 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05693 8185 8045 1496 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05692 2944 4470 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05691 2946 3033 2944 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05690 8185 1986 1664 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05689 1664 2926 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05688 3253 1802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05687 1664 1887 1802 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05686 1802 2698 1664 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05685 3026 4572 3027 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05684 3027 4051 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05683 3608 5483 3026 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05682 776 4572 775 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05681 775 4573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05680 1148 774 776 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05679 1548 6543 1549 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05678 1549 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05677 1553 2687 1548 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05676 7227 7328 7226 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05675 7226 7327 7326 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05674 8185 7329 7227 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05673 7325 7326 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05672 3040 4166 3039 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05671 3039 3759 3113 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05670 8185 3744 3040 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05669 3111 3113 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05668 3041 4424 3042 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05667 3042 3763 3125 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05666 8185 3744 3041 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05665 3123 3125 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05664 1244 1550 1245 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05663 1245 1361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05662 1243 1362 1244 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05661 1792 1553 1243 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05660 2440 2437 2442 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05659 2442 2441 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05658 2438 2693 2440 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05657 2439 2913 2438 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05656 6820 6821 6706 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05655 6706 7058 6820 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05654 8185 7053 6706 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05653 8185 1996 1581 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05652 1581 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05651 2233 1580 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05650 1581 1891 1580 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05649 1580 2926 1581 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05648 2577 6797 2578 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05647 2578 4575 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05646 2576 4167 2577 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05645 2723 4306 2576 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05644 5266 6172 5267 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05643 5267 6396 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05642 5264 6421 5266 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05641 5265 6921 5264 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05640 8185 2254 2031 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05639 2031 2252 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05638 2032 2031 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05637 4320 4583 4319 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05636 4319 5041 4320 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05635 8185 4317 4319 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05634 4318 4320 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05633 6513 6502 6505 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05632 6505 6503 6513 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05631 8185 6504 6505 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05630 6915 7305 6749 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05629 6749 7301 6915 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05628 8185 6914 6749 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05627 8185 2926 2920 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05626 8185 3171 2920 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05625 2920 3170 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05624 2919 2920 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05623 5900 6090 5636 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05622 5636 6089 5900 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05621 8185 6576 5636 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05620 4168 4167 4169 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05619 4169 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05618 4165 7353 4168 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05617 4166 6506 4165 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05616 7239 7884 7238 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05615 7238 7403 7402 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05614 8185 7883 7239 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05613 8179 7402 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05612 3715 3716 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05611 8185 7787 3715 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05610 3715 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05609 8185 8045 3715 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05608 3714 3715 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05607 8185 4405 4139 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05606 4139 4898 4138 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05605 4137 4138 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05604 8185 2924 1552 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05603 1552 1559 1551 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05602 1550 1551 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05601 8185 4572 2456 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05600 2456 2469 2455 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05599 2707 2455 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05598 8185 4574 2092 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05597 2092 6797 2218 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05596 2896 2218 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05595 8185 1043 1044 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05594 1044 5641 1045 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05593 1743 1045 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05592 6789 7280 6687 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05591 6687 6835 6789 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05590 8185 7025 6687 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05589 6788 6789 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05588 4018 7791 3916 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05587 3916 7788 4018 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05586 8185 6080 3916 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05585 5382 5380 5279 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05584 5279 5633 5382 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05583 8185 5817 5279 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05582 5379 5382 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05581 5423 5421 5302 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05580 5302 5633 5423 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05579 8185 7536 5302 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05578 5420 5423 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05577 8185 8184 5790 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05576 5790 8187 5975 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05575 5879 5975 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05574 45 1150 46 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05573 46 359 164 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05572 8185 3384 45 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05571 163 164 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05570 3739 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_05569 4143 3991 3739 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_05568 3738 3740 4143 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_05567 8185 3737 3738 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_05566 3738 4141 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_05565 5928 5929 5770 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05564 5770 6019 5928 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05563 8185 5927 5770 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05562 6102 5928 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05561 2251 2249 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05560 8185 2454 2251 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05559 4882 5041 4883 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05558 4883 5273 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05557 4881 5269 4882 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05556 5040 5043 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05555 5043 5042 4881 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05554 7323 7797 7171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05553 7171 7798 7323 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05552 8185 7585 7171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05551 2124 2269 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05550 2125 2270 2267 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05549 2123 2271 2264 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05548 8185 2262 2123 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05547 8185 3834 2271 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05546 2270 2271 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05545 8185 3193 2269 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05544 2267 2271 2124 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05543 2265 2267 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05542 8185 2265 2125 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05541 2264 2270 2265 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05540 2262 2264 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05539 8185 2264 2262 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05538 5206 5209 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05537 5208 5210 5207 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05536 5203 5211 5204 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05535 8185 5202 5203 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05534 8185 5864 5211 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05533 5210 5211 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05532 8185 5487 5209 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05531 5207 5211 5206 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05530 5205 5207 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05529 8185 5205 5208 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05528 5204 5210 5205 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05527 5202 5204 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05526 8185 5204 5202 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05525 4313 5265 4314 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05524 4314 4583 4313 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05523 8185 4312 4314 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05522 4311 4313 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05521 1895 5940 1896 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05520 1896 2262 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05519 1894 2964 1895 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05518 2469 2030 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05517 2030 2968 1894 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05516 2027 1897 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05515 8185 1898 2027 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05514 847 4573 848 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05513 848 4575 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05512 846 6609 847 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05511 1618 968 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05510 968 4302 846 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05509 3499 6797 3498 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05508 3498 3639 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05507 3497 6609 3499 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05506 3856 3640 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05505 3640 6293 3497 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05504 3132 3552 2999 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05503 2999 3141 3132 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05502 8185 3553 2999 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05501 3130 3132 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05500 3277 3276 3278 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05499 3278 3964 3277 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05498 8185 4503 3278 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05497 3275 3277 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05496 34 152 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05495 33 153 149 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05494 32 154 146 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05493 8185 532 32 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05492 8185 3834 154 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05491 153 154 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05490 8185 320 152 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05489 149 154 34 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05488 148 149 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05487 8185 148 33 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05486 146 153 148 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05485 532 146 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05484 8185 146 532 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05483 433 763 432 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05482 432 557 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05481 942 565 433 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05480 1536 4172 1534 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05479 1534 1782 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05478 1535 1539 1536 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05477 1542 4172 1540 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05476 1540 1538 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05475 1541 1539 1542 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05474 3061 3191 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05473 3193 3192 3061 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05472 4208 4021 3917 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05471 3917 7788 4208 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05470 8185 6541 3917 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05469 1465 5099 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05468 3958 1466 1465 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05467 3049 3150 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05466 3353 6363 3049 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05465 4950 7059 4838 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05464 4838 5406 4950 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05463 8185 6834 4838 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05462 4947 4950 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05461 4845 4974 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05460 4846 4975 4973 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05459 4844 4976 4969 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05458 8185 5180 4844 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05457 8185 5864 4976 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05456 4975 4976 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05455 8185 5181 4974 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05454 4973 4976 4845 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05453 4970 4973 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05452 8185 4970 4846 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05451 4969 4975 4970 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05450 5180 4969 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05449 8185 4969 5180 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05448 1485 1484 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05447 1482 1486 1483 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05446 1480 1487 1479 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05445 8185 5571 1480 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05444 8185 1951 1487 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05443 1486 1487 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05442 8185 1488 1484 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05441 1483 1487 1485 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05440 1481 1483 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05439 8185 1481 1482 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05438 1479 1486 1481 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05437 5571 1479 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05436 8185 1479 5571 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05435 4667 4668 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05434 4613 4615 4614 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05433 4611 4669 4665 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05432 8185 5108 4611 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05431 8185 8063 4669 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05430 4615 4669 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05429 8185 4666 4668 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05428 4614 4669 4667 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05427 4612 4614 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05426 8185 4612 4613 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05425 4665 4615 4612 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05424 5108 4665 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05423 8185 4665 5108 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05422 7749 7766 7658 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05421 7658 7747 7749 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05420 8185 7748 7658 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05419 5414 5413 5298 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05418 5298 5432 5414 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05417 8185 5436 5298 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05416 7695 7890 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05415 8175 7887 7695 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05414 7685 7878 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05413 7875 7874 7685 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05412 6748 6915 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05411 7399 6912 6748 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05410 6233 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05409 6627 6618 6233 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05408 3854 3867 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05407 3853 4292 3854 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05406 2630 4171 2061 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05405 2061 2167 2630 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05404 8185 2375 2061 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05403 3281 3284 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05402 3228 3283 3227 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05401 3225 3285 3279 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05400 8185 5563 3225 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05399 8185 3708 3285 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05398 3283 3285 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05397 8185 3282 3284 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05396 3227 3285 3281 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05395 3226 3227 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05394 8185 3226 3228 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05393 3279 3283 3226 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05392 5563 3279 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05391 8185 3279 5563 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05390 8185 7343 7032 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05389 7032 7053 7031 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05388 7339 7031 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05387 6220 7356 6219 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05386 6219 6311 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05385 6218 7051 6220 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05384 7034 6349 6218 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05383 6232 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05382 6897 6883 6232 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05381 5358 6415 5357 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05380 5357 5500 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05379 5501 6412 5358 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05378 1574 5654 1573 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05377 1573 7026 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05376 1806 7353 1574 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05375 6752 7408 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05374 7149 8184 6752 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05373 6113 6838 6343 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05372 8185 6343 6590 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05371 8185 6838 6346 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05370 6114 6344 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05369 6343 6346 6114 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05368 8185 6341 6113 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05367 6590 6343 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05366 6589 6864 6592 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05365 8185 6592 6597 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05364 8185 6864 6593 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05363 6591 6590 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05362 6592 6593 6591 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05361 8185 6588 6589 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05360 6597 6592 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05359 3503 3660 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05358 3661 4074 3503 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05357 8185 6090 4948 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05356 4837 4948 4946 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05355 8185 7343 4837 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05354 4945 4946 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05353 8185 4946 4945 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05352 4836 5147 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05351 4943 5148 4836 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05350 8185 7955 4943 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05349 4942 4943 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05348 8185 3553 2343 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05347 2343 3097 2345 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05346 2344 2345 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05345 8185 3229 2995 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05344 2995 3316 3117 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05343 3559 3117 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05342 3762 4172 3764 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05341 3764 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05340 3763 7863 3762 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05339 13 903 94 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05338 8185 94 91 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05337 8185 903 95 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05336 14 3532 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05335 94 95 14 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05334 8185 268 13 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05333 91 94 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05332 6695 7026 6694 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05331 6694 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05330 6693 6796 6695 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05329 7012 8000 6693 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05328 1047 1476 1046 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05327 1046 1477 1047 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05326 8185 8045 1046 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05325 770 4306 771 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05324 771 6609 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05323 1891 5447 770 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05322 5968 7893 5786 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05321 5786 7408 5968 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05320 8185 8184 5786 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05319 5271 6396 5270 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05318 5270 5875 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05317 5268 6172 5271 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05316 5269 6672 5268 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05315 6569 6838 6568 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05314 8185 6568 6588 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05313 8185 6838 6571 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05312 6570 6823 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05311 6568 6571 6570 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05310 8185 6567 6569 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05309 6588 6568 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05308 3838 4061 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05307 3867 3841 3838 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05306 8185 4280 3867 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05305 1812 2926 1667 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05304 1667 1996 1812 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05303 8185 1813 1667 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05302 2239 1812 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05301 2431 4293 2429 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05300 2429 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05299 2430 2968 2431 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05298 2000 5483 2001 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05297 2001 4293 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05296 1999 5940 2000 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05295 7494 7729 7495 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05294 7495 7734 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05293 7493 7738 7494 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05292 7742 7730 7493 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05291 3295 4178 3535 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05290 8185 3535 3532 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05289 8185 4178 3536 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05288 3296 4403 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05287 3535 3536 3296 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05286 8185 7528 3295 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05285 3532 3535 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05284 6527 7026 6528 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05283 6528 6543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05282 6526 6544 6527 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05281 6794 8021 6526 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05280 3478 7356 3479 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05279 3479 3639 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05278 3477 6609 3478 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05277 3618 6293 3477 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05276 6522 6797 6523 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05275 6523 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05274 6521 6796 6522 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05273 7006 6520 6521 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05272 3365 5168 3364 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05271 3364 3608 3366 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05270 8185 3373 3365 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05269 3610 3366 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05268 8185 3556 1639 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05267 1724 1719 1637 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05266 1722 2813 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_05265 1637 1721 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05264 8185 3556 1721 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_05263 2589 1724 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_05262 1639 1727 1638 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05261 1638 2813 1724 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05260 1724 1722 1640 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05259 1640 2610 1639 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_05258 3892 3985 4149 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05257 8185 3986 3892 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05256 3891 4143 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05255 4149 3983 3891 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05254 8185 4143 3985 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05253 3983 3986 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05252 262 903 264 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05251 8185 264 261 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05250 8185 903 265 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05249 263 3978 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05248 264 265 263 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05247 8185 498 262 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05246 261 264 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05245 4713 7314 6850 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05244 8185 7314 4715 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05243 4716 4714 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05242 6850 4715 4716 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05241 8185 4712 4713 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05240 8185 5606 5123 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05239 5123 5121 5122 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05238 5120 5122 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05237 8185 6576 5768 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05236 5768 6127 5920 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05235 5846 5920 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05234 8185 5900 5755 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05233 5755 6288 5899 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05232 5828 5899 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05231 7762 7761 7660 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05230 7660 7760 7762 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05229 8185 7979 7660 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05228 7759 7762 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05227 5100 6524 5101 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05226 5101 5406 5100 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05225 8185 5124 5101 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05224 5099 5100 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05223 243 246 1287 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05222 8185 1711 243 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05221 245 1924 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05220 1287 244 245 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05219 8185 1924 246 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05218 244 1711 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05217 3971 6541 3888 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05216 8185 8064 3973 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05215 3888 3973 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05214 8185 3078 645 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05213 645 2315 646 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05212 2806 646 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05211 8185 4572 2573 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05210 2573 2719 2717 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05209 2937 2717 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05208 8185 2235 1670 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05207 1670 2027 1814 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05206 1817 1814 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05205 3765 6484 3766 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05204 8185 8064 3767 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05203 3766 3767 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05202 6045 6050 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05201 6044 6262 6045 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05200 8185 6274 6044 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05199 6043 6044 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05198 6781 6500 6501 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05197 6501 6783 6781 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05196 8185 7314 6501 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05195 4387 5938 4386 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05194 4386 5453 4486 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05193 8185 5606 4387 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05192 4402 4486 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05191 8185 7891 6634 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05190 6634 7881 6633 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05189 6632 6633 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05188 5812 7893 5813 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05187 5813 8187 5972 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05186 8185 7883 5812 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05185 5875 5972 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05184 8185 7130 5371 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05183 5371 7633 5510 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05182 6912 5510 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05181 819 5483 818 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05180 818 4302 953 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05179 8185 5940 819 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05178 1133 953 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05177 8185 1546 5620 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05176 5620 1547 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05175 8185 1545 5620 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05174 8185 6334 6224 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05173 6224 7788 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05172 6329 6331 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05171 6224 6340 6331 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05170 6331 6332 6224 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05169 5214 5695 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05168 5213 5869 5214 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05167 8185 5212 5213 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05166 7863 7591 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05165 8122 8058 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05164 3823 4302 3822 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05163 3822 6609 3824 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05162 8185 5654 3823 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05161 7788 3824 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_05160 3877 2950 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05159 8185 2951 3877 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05158 2709 5492 2570 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05157 2571 4295 2709 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05156 2570 4790 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05155 2705 2709 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05154 8185 2707 2571 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05153 2571 2706 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_05152 1153 1543 1155 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05151 1155 1154 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05150 1151 1559 1153 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05149 1150 1152 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_05148 1152 1806 1151 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05147 804 873 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05146 803 874 871 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05145 802 875 868 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05144 8185 1048 802 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05143 8185 1951 875 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05142 874 875 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05141 8185 890 873 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05140 871 875 804 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05139 869 871 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05138 8185 869 803 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05137 868 874 869 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05136 1048 868 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05135 8185 868 1048 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05134 7366 7791 7194 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05133 7194 7788 7366 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05132 8185 8097 7194 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05131 7368 7366 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05130 7112 7379 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05129 8185 342 336 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05128 336 343 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05127 1110 335 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05126 336 334 335 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05125 335 354 336 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05124 4158 4498 4159 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05123 4159 4157 4158 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05122 8185 4155 4159 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05121 4156 4158 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05120 3385 3386 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05119 3243 3387 3242 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05118 3240 3388 3382 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05117 8185 3384 3240 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05116 8185 3834 3388 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05115 3387 3388 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05114 8185 4757 3386 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05113 3242 3388 3385 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05112 3241 3242 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05111 8185 3241 3243 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05110 3382 3387 3241 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05109 3384 3382 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05108 8185 3382 3384 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05107 5303 6480 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05106 5424 5603 5303 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05105 3046 3146 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05104 3141 4007 3046 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05103 20 111 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05102 19 112 110 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05101 18 113 106 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05100 8185 703 18 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05099 8185 1951 113 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05098 112 113 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05097 8185 697 111 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05096 110 113 20 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05095 107 110 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05094 8185 107 19 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05093 106 112 107 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05092 703 106 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05091 8185 106 703 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05090 1032 1036 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05089 1034 1035 1033 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05088 1029 1037 1030 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05087 8185 6267 1029 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05086 8185 3708 1037 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05085 1035 1037 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05084 8185 6085 1036 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05083 1033 1037 1032 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05082 1031 1033 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05081 8185 1031 1034 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05080 1030 1035 1031 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05079 6267 1030 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05078 8185 1030 6267 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05077 5659 6358 5661 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05076 8185 5661 5658 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05075 8185 6358 5662 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05074 5660 6076 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05073 5661 5662 5660 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05072 8185 6142 5659 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05071 5658 5661 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05070 2069 4693 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05069 2182 2181 2069 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05068 2564 3158 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05067 2702 3857 2564 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05066 3043 3768 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05065 3129 3128 3043 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05064 7212 7393 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05063 7211 7389 7392 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05062 7210 7390 7388 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05061 8185 7604 7210 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05060 8185 8166 7390 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05059 7389 7390 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05058 8185 7603 7393 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05057 7392 7390 7212 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05056 7391 7392 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05055 8185 7391 7211 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05054 7388 7389 7391 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05053 7604 7388 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05052 8185 7388 7604 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05051 8185 1372 1137 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05050 1137 3608 1138 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05049 1359 1138 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05048 4272 7871 4273 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05047 8185 4273 4271 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05046 8185 7871 4275 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05045 4274 4788 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05044 4273 4275 4274 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05043 8185 4270 4272 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_05042 4271 4273 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05041 5117 5606 5119 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05040 5119 5121 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05039 5118 6549 5117 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05038 4796 7887 4797 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05037 4797 6421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05036 4795 5740 4796 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05035 8185 6667 6187 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05034 6187 6188 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05033 6185 6186 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05032 6187 7299 6186 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05031 6186 6189 6187 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_05030 3915 6089 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05029 4202 4029 3915 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05028 8185 6090 4202 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05027 3012 5168 3011 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05026 3011 3608 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05025 3780 3373 3012 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05024 8185 5168 5170 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05023 5170 5169 5171 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05022 6835 5171 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05021 6966 6970 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05020 6968 6969 6967 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05019 6963 6971 6964 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05018 8185 7247 6963 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05017 8185 8063 6971 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05016 6969 6971 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_05015 8185 7241 6970 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_05014 6967 6971 6966 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05013 6965 6967 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05012 8185 6965 6968 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05011 6964 6969 6965 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_05010 7247 6964 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05009 8185 6964 7247 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05008 8185 7343 7045 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05007 7045 7062 7046 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05006 7543 7046 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05005 5079 6477 5080 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05004 5080 5078 5079 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05003 8185 7957 5080 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05002 5077 5079 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_05001 4884 6921 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_05000 5044 7130 4884 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04999 3487 7356 3486 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04998 3486 3826 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04997 3485 4306 3487 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04996 3623 5942 3485 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04995 3935 6311 3936 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04994 3936 4047 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04993 3934 4573 3935 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04992 4048 6293 3934 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04991 8185 1799 381 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04990 380 381 379 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04989 8185 2492 380 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04988 378 379 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04987 8185 379 378 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04986 8185 7343 2451 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04985 2451 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04984 2448 2452 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04983 2451 4517 2452 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04982 2452 2926 2451 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04981 6302 6090 6091 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04980 6091 6089 6302 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04979 8185 6823 6091 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04978 8185 7512 7510 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04977 7510 7508 7509 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04976 7753 7509 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04975 3899 4574 3900 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04974 3900 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04973 3898 6293 3899 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04972 3990 6775 3898 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04971 1948 3114 2164 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04970 8185 2164 2166 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04969 8185 3114 2162 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04968 1950 3348 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04967 2164 2162 1950 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04966 8185 3315 1948 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04965 2166 2164 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04964 8185 7343 5750 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04963 5750 5896 5895 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04962 5825 5895 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04961 2909 3378 2908 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04960 2908 4517 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04959 2907 3379 2909 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04958 2906 5169 2907 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04957 4372 7871 4576 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04956 8185 4576 4570 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04955 8185 7871 4466 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04954 4373 6648 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04953 4576 4466 4373 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04952 8185 4734 4372 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04951 4570 4576 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04950 5487 6629 5342 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04949 5342 5494 5487 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04948 8185 5486 5342 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04947 8185 2492 374 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04946 373 374 372 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04945 8185 1799 373 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04944 375 372 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04943 8185 372 375 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04942 8185 4302 3013 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04941 3013 5624 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04940 7797 3152 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04939 3013 3370 3152 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04938 3152 3371 3013 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_04937 825 1154 826 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04936 826 4228 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04935 824 5147 825 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04934 955 1543 824 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04933 7087 7867 7088 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04932 8185 7088 7398 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04931 8185 7867 7090 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04930 7089 7528 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04929 7088 7090 7089 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04928 8185 7572 7087 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04927 7398 7088 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04926 4204 4705 4205 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04925 4205 4203 4204 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04924 8185 4202 4205 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04923 4206 4204 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04922 2420 2421 2419 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04921 2419 2430 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04920 2418 4203 2420 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04919 5406 2417 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04918 2417 2924 2418 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04917 4820 4902 4821 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04916 4821 4901 4903 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04915 8185 5606 4820 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04914 4900 4903 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04913 3953 5483 3952 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04912 3952 5447 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04911 3951 7051 3953 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04910 4583 4075 3951 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04909 8185 4298 4300 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04908 4300 4473 4301 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04907 4299 4301 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04906 8185 4956 4343 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04905 4343 5399 4516 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04904 4437 4516 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04903 679 1115 681 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04902 681 1114 680 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04901 680 1063 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04900 678 676 681 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04899 8185 1110 678 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04898 8185 677 679 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04897 1477 681 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04896 2158 2156 2056 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04895 2056 2822 2158 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04894 8185 3315 2056 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04893 2155 2158 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04892 2177 1964 1961 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04891 1961 1965 2177 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04890 8185 1962 1961 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04889 3326 3323 3577 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04888 8185 3567 3326 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04887 3325 3570 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04886 3577 3324 3325 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04885 8185 3570 3323 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04884 3324 3567 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04883 6279 6489 6198 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04882 8185 7500 6277 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04881 6198 6277 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04880 8185 5606 5282 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04879 5282 5384 5385 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04878 5390 5385 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04877 1264 7026 1263 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04876 1263 4575 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04875 1262 4572 1264 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04874 1377 1378 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04873 1378 5447 1262 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04872 3248 5648 3247 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04871 3247 6543 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04870 3246 6544 3248 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04869 3390 3389 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04868 3389 3857 3246 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04867 3367 6609 3368 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04866 3368 4068 3369 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04865 8185 4293 3367 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04864 4021 3369 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04863 2974 2975 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04862 2973 2976 2972 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04861 2969 2977 2970 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04860 8185 2968 2969 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04859 8185 3834 2977 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04858 2976 2977 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04857 8185 3197 2975 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04856 2972 2977 2974 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04855 2971 2972 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04854 8185 2971 2973 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04853 2970 2976 2971 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04852 2968 2970 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04851 8185 2970 2968 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04850 8185 8064 467 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04849 389 467 466 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04848 8185 3077 389 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04847 1909 466 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04846 8185 466 1909 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04845 6815 7779 6705 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04844 6705 7778 6815 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04843 8185 7349 6705 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04842 6816 6815 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04841 2953 4468 2956 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04840 2956 2955 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04839 2954 2958 2953 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04838 3186 2952 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04837 2952 2957 2954 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04836 8185 2696 2917 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04835 2917 2904 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04834 8185 2695 2917 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04833 8185 2919 3167 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04832 3167 2917 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04831 8185 3251 3167 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04830 8185 3644 3189 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04829 3035 3189 3188 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04828 8185 3187 3035 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04827 3191 3188 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04826 8185 3188 3191 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04825 2476 2723 2478 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04824 2478 2722 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04823 2474 2481 2476 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04822 2471 2475 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04821 2475 2473 2474 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04820 7100 7103 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04819 7099 7102 7101 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04818 7096 7105 7097 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04817 8185 7095 7096 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04816 8185 8166 7105 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04815 7102 7105 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04814 8185 7108 7103 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04813 7101 7105 7100 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04812 7098 7101 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04811 8185 7098 7099 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04810 7097 7102 7098 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04809 7095 7097 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04808 8185 7097 7095 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04807 4941 4939 4835 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04806 4835 6294 4941 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04805 8185 5144 4835 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04804 5428 4941 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04803 1890 2216 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04802 8185 2005 1890 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04801 1890 1889 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04800 8185 2439 1890 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04799 2436 7353 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04798 2441 3371 2436 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04797 2435 4302 2441 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04796 8185 2682 2435 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04795 2434 2896 2441 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04794 8185 4306 2434 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04793 6836 7591 6710 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04792 6710 6835 6836 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04791 8185 7062 6710 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04790 6834 6836 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04789 1625 1626 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04788 1624 1627 1623 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04787 1620 1628 1621 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04786 8185 1799 1620 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04785 8185 3834 1628 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04784 1627 1628 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04783 8185 2961 1626 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04782 1623 1628 1625 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04781 1622 1623 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04780 8185 1622 1624 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04779 1621 1627 1622 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04778 1799 1621 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04777 8185 1621 1799 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04776 1656 1770 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04775 1655 1773 1768 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04774 1654 1774 1766 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04773 8185 5435 1654 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04772 8185 1772 1774 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04771 1773 1774 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04770 8185 1974 1770 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04769 1768 1774 1656 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04768 1767 1768 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04767 8185 1767 1655 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04766 1766 1773 1767 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04765 5435 1766 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04764 8185 1766 5435 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04763 2326 2328 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04762 2323 2327 2325 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04761 2321 2329 2322 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04760 8185 6292 2321 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04759 8185 3708 2329 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04758 2327 2329 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04757 8185 4641 2328 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04756 2325 2329 2326 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04755 2324 2325 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04754 8185 2324 2323 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04753 2322 2327 2324 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04752 6292 2322 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04751 8185 2322 6292 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04750 773 1543 772 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04749 772 778 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04748 946 1157 773 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04747 3375 5654 3374 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04746 3374 5648 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04745 3373 7051 3375 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04744 4581 4583 4385 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04743 4385 5038 4581 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04742 8185 4582 4385 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04741 4477 4581 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04740 4175 4172 4174 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04739 4174 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04738 4511 7777 4175 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04737 811 1123 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04736 923 1110 811 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04735 7070 7263 7069 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_04734 7071 7550 7070 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_04733 7069 7264 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_04732 7068 7070 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_04731 8185 7548 7071 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_04730 7071 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_04729 437 5654 436 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04728 436 4293 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04727 1157 5483 437 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04726 3245 3390 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04725 3244 6598 3245 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04724 8185 3583 3585 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04723 3460 3585 3584 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04722 8185 3776 3460 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04721 3582 3584 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04720 8185 3584 3582 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04719 5293 7247 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04718 5399 6285 5293 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04717 5292 6286 5399 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04716 8185 6506 5292 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04715 5291 6801 5399 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04714 8185 6284 5291 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04713 3430 3520 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04712 3431 3521 3517 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04711 3429 3522 3514 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04710 8185 5387 3429 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04709 8185 3708 3522 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04708 3521 3522 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04707 8185 3519 3520 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04706 3517 3522 3430 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04705 3515 3517 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04704 8185 3515 3431 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04703 3514 3521 3515 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04702 5387 3514 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04701 8185 3514 5387 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04700 6698 7356 6699 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04699 6699 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04698 6697 7353 6698 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04697 7333 6801 6697 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04696 8185 5618 5621 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04695 5621 5620 5622 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04694 5619 5622 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04693 5719 6900 5717 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04692 5717 8187 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04691 5718 7883 5719 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04690 2465 2469 2464 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04689 2464 4575 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04688 2462 4302 2465 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04687 8185 2951 2479 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04686 2479 2950 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04685 2477 2479 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04684 1532 5148 1533 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04683 1533 2203 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04682 2202 1986 1532 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04681 7317 7955 7167 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04680 7167 7747 7317 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04679 8185 7319 7167 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04678 7489 7317 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04677 8185 3556 2052 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04676 2149 2144 2049 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04675 2147 2813 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_04674 2049 2145 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04673 8185 3556 2145 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_04672 2143 2149 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_04671 2052 2337 2050 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04670 2050 2813 2149 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04669 2149 2147 2051 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04668 2051 2340 2052 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04667 8185 6359 4750 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04666 4992 7612 4746 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04665 4990 4997 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_04664 4746 4988 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04663 8185 6359 4988 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_04662 4987 4992 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_04661 4750 5202 4748 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04660 4748 4997 4992 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04659 4992 4990 4747 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04658 4747 7056 4750 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_04657 3889 4178 3979 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04656 8185 3979 3978 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04655 8185 4178 3982 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04654 3890 5391 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04653 3979 3982 3890 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04652 8185 7585 3889 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04651 3978 3979 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04650 7027 7026 7028 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04649 7028 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04648 7024 7051 7027 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04647 7025 8040 7024 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04646 4140 4712 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04645 4507 7314 4140 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04644 4284 7354 4285 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04643 4285 4575 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04642 4283 4306 4284 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04641 4286 5654 4283 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04640 4866 6921 4865 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04639 4865 6636 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04638 4864 5868 4866 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04637 5031 7130 4864 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04636 4793 4790 4794 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04635 4794 6421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04634 4791 7887 4793 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04633 4792 7149 4791 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04632 4142 4146 4497 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04631 8185 4141 4142 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04630 4145 4143 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04629 4497 4144 4145 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04628 8185 4143 4146 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04627 4144 4141 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04626 2841 3759 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04625 2842 4166 2841 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04624 8185 4510 2842 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04623 2840 2842 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04622 428 903 550 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04621 8185 550 751 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04620 8185 903 465 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04619 429 4012 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04618 550 465 429 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04617 8185 1116 428 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04616 751 550 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04615 3913 5148 4014 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04614 8185 4014 4012 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04613 8185 5148 4016 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04612 3914 7349 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04611 4014 4016 3914 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04610 8185 6541 3913 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04609 4012 4014 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04608 702 903 901 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04607 8185 901 899 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04606 8185 903 905 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04605 704 4160 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04604 901 905 704 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04603 8185 900 702 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04602 899 901 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04601 4161 4178 4162 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04600 8185 4162 4160 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04599 8185 4178 4164 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04598 4163 4414 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04597 4162 4164 4163 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04596 8185 7777 4161 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04595 4160 4162 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04594 8185 4428 4185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04593 4185 5837 4187 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04592 4184 4187 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04591 5412 5413 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04590 8185 7787 5412 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04589 5412 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04588 8185 8045 5412 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04587 5408 5412 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04586 6989 7957 6988 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04585 8185 7957 6991 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04584 6990 6992 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04583 6988 6991 6990 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04582 8185 6987 6989 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04581 1610 4068 1609 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04580 1609 4295 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04579 1608 7026 1610 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04578 1611 6796 1608 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04577 3649 3851 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04576 8185 3853 3649 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04575 3649 3645 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04574 8185 3651 3649 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04573 3644 3649 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04572 8185 2466 2468 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04571 8185 2705 2468 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04570 2468 2467 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04569 2962 2468 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04568 7512 7797 7511 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04567 7511 7798 7512 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04566 8185 7549 7511 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04565 800 866 865 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04564 8185 2136 800 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04563 801 1924 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04562 865 863 801 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04561 8185 1924 866 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04560 863 2136 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04559 8185 965 966 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04558 6802 966 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04557 8185 966 6802 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04556 8185 966 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04555 8144 966 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04554 8185 965 784 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04553 6311 784 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04552 8185 784 6311 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04551 8185 784 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04550 8144 784 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04549 8185 574 572 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04548 965 572 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04547 8185 572 965 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04546 8185 572 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04545 8144 572 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04544 8185 7314 6275 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04543 6197 6275 6276 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04542 8185 6273 6197 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04541 6274 6276 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04540 8185 6276 6274 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04539 8185 1799 779 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04538 779 2492 780 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04537 2718 780 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04536 4780 5720 4781 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04535 4781 4782 4780 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04534 8185 7352 4781 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04533 4779 4780 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04532 8185 4792 3848 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04531 3848 3847 3849 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04530 3850 3849 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04529 8185 7885 7216 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04528 7216 7877 7396 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04527 7299 7396 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04526 8185 3860 3505 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04525 3505 3868 3666 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04524 3665 3666 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04523 8185 5838 5601 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04522 5601 6062 5602 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04521 5600 5602 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04520 8185 7645 6922 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04519 6921 6922 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04518 8185 6922 6921 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04517 8185 6922 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04516 8144 6922 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04515 8185 7645 6673 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04514 6672 6673 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04513 8185 6673 6672 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04512 8185 6673 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04511 8144 6673 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04510 8185 7646 7647 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04509 7645 7647 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04508 8185 7647 7645 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04507 8185 7647 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04506 8144 7647 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04505 7155 7881 7156 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04504 7156 7403 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04503 7154 7884 7155 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04502 7405 7153 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04501 7153 8184 7154 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04500 7144 7888 7143 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04499 7143 7643 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04498 7142 8187 7144 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04497 7140 7141 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04496 7141 7883 7142 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04495 2414 2678 2415 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04494 2415 4018 2416 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04493 8185 2412 2414 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04492 2413 2416 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04491 8185 5908 2903 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04490 2903 2901 2902 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04489 2912 2902 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04488 4732 4955 4733 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04487 4733 4730 4732 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04486 8185 4731 4733 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04485 5680 4732 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04484 444 4228 445 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04483 445 760 556 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04482 8185 1891 444 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04481 559 556 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04480 5396 6793 5290 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04479 5290 5406 5396 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04478 8185 6517 5290 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04477 5395 5396 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04476 2461 2469 2460 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04475 2460 4575 2463 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04474 8185 4302 2461 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04473 2710 2463 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04472 7119 7604 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04471 8137 8147 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04470 7596 8125 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04469 5704 6629 5705 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04468 5705 5710 5704 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04467 8185 5862 5705 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04466 7858 8119 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04465 5025 5015 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04464 4635 4558 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04463 3391 4270 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04462 4251 3384 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04461 5000 5485 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04460 1818 2039 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04459 8185 1893 1818 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04458 2154 2156 2055 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04457 2055 2822 2154 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04456 8185 3315 2055 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04455 2066 4003 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04454 2379 2177 2066 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04453 3329 3552 3328 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04452 3328 3327 3329 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04451 8185 3553 3328 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04450 3569 3329 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04449 3752 3750 3753 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04448 3753 3751 3752 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04447 8185 8064 3753 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04446 4326 6867 4666 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04445 8185 6867 4491 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04444 4327 4492 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04443 4666 4491 4327 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04442 8185 4901 4326 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04441 1023 1024 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04440 1021 1026 1022 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04439 1018 1025 1019 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04438 8185 1043 1018 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04437 8185 3708 1025 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04436 1026 1025 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04435 8185 1038 1024 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04434 1022 1025 1023 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04433 1020 1022 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04432 8185 1020 1021 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04431 1019 1026 1020 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04430 1043 1019 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04429 8185 1019 1043 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04428 3833 3832 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04427 3830 3835 3831 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04426 3827 3836 3828 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04425 8185 4270 3827 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04424 8185 3834 3836 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04423 3835 3836 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04422 8185 4271 3832 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04421 3831 3836 3833 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04420 3829 3831 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04419 8185 3829 3830 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04418 3828 3835 3829 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04417 4270 3828 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04416 8185 3828 4270 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04415 7186 7352 7187 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04414 7187 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04413 7340 8086 7186 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04412 5365 7405 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04411 5507 7633 5365 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04410 1353 2492 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04409 7963 7966 7964 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04408 7964 7962 7963 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04407 8185 7960 7964 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04406 1471 1943 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04405 1470 2154 1471 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04404 8185 2616 1470 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04403 1732 1470 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04402 2846 3570 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04401 3118 2845 2846 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04400 1240 1356 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04399 1547 1553 1240 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04398 823 957 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04397 1546 4540 823 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04396 1544 5169 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04395 1545 1543 1544 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04394 5623 7883 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04393 5629 7352 5623 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04392 945 943 816 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04391 816 942 945 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04390 8185 1119 816 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04389 1120 945 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04388 6098 6325 6327 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04387 8185 6327 6563 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04386 8185 6325 6328 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04385 6099 6329 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04384 6327 6328 6099 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04383 8185 6567 6098 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04382 6563 6327 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04381 4861 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04380 5026 5025 4861 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04379 4863 5242 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04378 5030 5872 4863 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04377 1028 4651 1027 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04376 1027 5377 1028 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04375 8185 3968 1027 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04374 4658 1028 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04373 7775 7791 7662 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04372 7662 7788 7775 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04371 8185 8000 7662 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04370 7774 7775 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04369 2378 2847 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04368 2382 3229 2378 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04367 6039 6040 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04366 6009 6011 6010 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04365 6007 6041 6038 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04364 8185 6273 6007 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04363 8185 8063 6041 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04362 6011 6041 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04361 8185 6043 6040 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04360 6010 6041 6039 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04359 6008 6010 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04358 8185 6008 6009 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04357 6038 6011 6008 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04356 6273 6038 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04355 8185 6038 6273 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04354 8185 7252 7023 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04353 7023 7033 7022 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04352 7517 7022 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04351 6109 6359 6336 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04350 8185 6336 6334 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04349 8185 6359 6339 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04348 6110 7863 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04347 6336 6339 6110 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04346 8185 6335 6109 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04345 6334 6336 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04344 3238 3608 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04343 7791 5168 3238 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04342 1239 1365 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04341 2889 1550 1239 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04340 2101 2232 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04339 2712 2233 2101 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04338 8185 7343 7015 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04337 7015 7025 7016 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04336 7329 7016 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04335 8185 7957 7746 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04334 7657 7746 7745 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04333 8185 7979 7657 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04332 7744 7745 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04331 8185 7745 7744 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04330 7173 7352 7174 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04329 7174 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04328 7250 8000 7173 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04327 8155 8154 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04326 8151 8157 8152 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04325 8149 8158 8148 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04324 8185 8147 8149 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04323 8185 8166 8158 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04322 8157 8158 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04321 8185 8153 8154 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04320 8152 8158 8155 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04319 8150 8152 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04318 8185 8150 8151 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04317 8148 8157 8150 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04316 8147 8148 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04315 8185 8148 8147 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04314 4126 4125 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04313 4123 4127 4124 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04312 4121 4128 4120 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04311 8185 7752 4121 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04310 8185 8063 4128 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04309 4127 4128 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04308 8185 7492 4125 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04307 4124 4128 4126 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04306 4122 4124 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04305 8185 4122 4123 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04304 4120 4127 4122 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04303 7752 4120 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04302 8185 4120 7752 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04301 8185 7343 5283 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04300 5283 5388 5386 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04299 5553 5386 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04298 947 1798 757 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04297 757 7548 947 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04296 8185 6363 757 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04295 4775 7871 4776 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04294 8185 4776 5232 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04293 8185 7871 4777 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04292 4778 7405 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04291 4776 4777 4778 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04290 8185 5227 4775 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04289 5232 4776 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04288 4772 7871 4771 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04287 8185 4771 4769 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04286 8185 7871 4773 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04285 4774 5241 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04284 4771 4773 4774 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04283 8185 4770 4772 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04282 4769 4771 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04281 4749 4997 4751 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04280 4751 5668 4749 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04279 8185 4998 4751 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04278 7628 7888 7629 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04277 7629 7643 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04276 7626 8187 7628 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04275 7627 7883 7626 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04274 6136 6138 6135 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04273 6135 6133 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04272 6134 6161 6136 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04271 6132 7887 6134 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04270 5280 5938 5281 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04269 5281 5453 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04268 5383 5606 5280 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04267 3078 7787 2979 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04266 2979 5907 3078 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04265 8185 6520 2979 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04264 7072 7867 7074 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04263 8185 7074 7403 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04262 8185 7867 7077 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04261 7075 7073 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04260 7074 7077 7075 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04259 8185 7270 7072 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04258 7403 7074 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04257 7583 7867 7584 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04256 8185 7584 7881 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04255 8185 7867 7588 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04254 7586 7585 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04253 7584 7588 7586 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04252 8185 7845 7583 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04251 7881 7584 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04250 5370 6920 5369 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04249 5369 6421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04248 5509 5740 5370 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04247 2989 3730 2988 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04246 2988 3735 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04245 2987 3586 2989 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04244 3097 3581 2987 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04243 5557 5559 5919 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04242 8185 6524 5557 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04241 5556 5558 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04240 5919 5555 5556 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04239 8185 5558 5559 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04238 5555 6524 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04237 5775 6293 5776 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04236 5776 5942 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04235 5774 5940 5775 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04234 5937 7314 5774 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04233 1995 6796 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04232 3797 2210 1995 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04231 1993 1992 3797 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04230 8185 4067 1993 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04229 1991 4293 3797 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04228 8185 2469 1991 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04227 7200 7867 7376 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04226 8185 7376 7892 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04225 8185 7867 7282 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04224 7201 7280 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04223 7376 7282 7201 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04222 8185 7581 7200 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_04221 7892 7376 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04220 4296 6543 4297 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04219 4297 4295 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04218 4294 4293 4296 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04217 4312 5648 4294 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04216 7008 7006 7010 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04215 7010 7017 7009 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04214 8185 7007 7008 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04213 7321 7009 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04212 6261 6262 6192 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04211 6192 6265 6261 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04210 8185 6260 6192 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04209 8185 5245 5243 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04208 5243 5249 5244 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04207 5242 5244 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04206 8185 6654 6657 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04205 6657 8179 6656 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04204 6655 6656 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04203 8185 6883 5177 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04202 5177 5445 5179 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04201 5176 5179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04200 7786 7955 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04199 8185 7787 7786 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04198 7786 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04197 8185 8045 7786 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04196 8025 7786 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04195 2482 5447 2483 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04194 2483 4067 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04193 2480 5942 2482 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04192 2481 4075 2480 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04191 2112 5648 2111 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04190 2111 4295 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04189 2110 4067 2112 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04188 2473 5447 2110 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04187 4688 6821 4689 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04186 4689 5406 4688 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04185 8185 6809 4689 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04184 6670 8187 6259 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04183 6259 7408 6670 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04182 8185 7891 6259 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04181 4827 4928 4925 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04180 8185 5118 4827 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04179 4828 4924 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04178 4925 4923 4828 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04177 8185 4924 4928 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04176 4923 5118 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04175 8185 7026 1661 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04174 1661 4573 1787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04173 1992 1787 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04172 1301 1743 1208 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04171 1208 1744 1301 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04170 8185 1962 1208 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04169 7796 7797 7666 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04168 7666 7798 7796 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04167 8185 7863 7666 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04166 5286 5393 5391 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04165 8185 7020 5286 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04164 5287 5390 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04163 5391 5389 5287 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04162 8185 5390 5393 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04161 5389 7020 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04160 8185 4790 2933 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04159 2933 5496 2934 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04158 2932 2934 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04157 8185 3857 2567 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04156 2567 2922 2704 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04155 2703 2704 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04154 1234 5148 1233 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04153 1233 2203 1350 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04152 8185 1986 1234 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04151 1355 1350 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04150 5679 6293 5678 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04149 5678 5942 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04148 5677 5940 5679 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04147 6138 5676 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04146 5676 7314 5677 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04145 6036 7884 6037 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04144 6037 7398 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04143 6035 6893 6036 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04142 6176 6174 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04141 6174 7891 6035 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04140 5324 5942 5323 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04139 5323 5447 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04138 5322 6796 5324 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04137 5445 5448 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04136 5448 6358 5322 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04135 3942 4068 3943 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04134 3943 6311 4063 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04133 8185 6293 3942 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04132 4061 4063 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04131 1275 2718 1274 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04130 1274 2719 1387 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04129 8185 3857 1275 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04128 1615 1387 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04127 5806 6900 5805 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04126 5805 8187 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04125 5804 7408 5806 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04124 5867 5965 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04123 5965 7891 5804 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04122 2333 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_04121 2591 2334 2333 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_04120 2332 2344 2591 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_04119 8185 3737 2332 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_04118 2332 2589 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_04117 4849 4984 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04116 4848 4985 4982 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04115 4847 4986 4978 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04114 8185 7867 4847 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04113 8185 5864 4986 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04112 4985 4986 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04111 8185 4983 4984 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04110 4982 4986 4849 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04109 4979 4982 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04108 8185 4979 4848 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04107 4978 4985 4979 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04106 7867 4978 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04105 8185 4978 7867 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04104 1171 6311 1174 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04103 1174 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04102 1172 4573 1171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04101 1169 1170 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04100 1170 4067 1172 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04099 5348 6900 5350 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04098 5350 8187 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04097 5349 6893 5348 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04096 5496 5497 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_04095 5497 7883 5349 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04094 5320 5942 5321 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04093 5321 5447 5446 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04092 8185 7353 5320 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04091 5916 5446 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_04090 2453 4517 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04089 8185 2698 2453 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04088 2453 5147 2454 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04087 2454 2926 2453 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04086 7967 7965 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04085 7966 8064 7967 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04084 2371 2174 2064 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04083 2064 4183 2371 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04082 8185 2365 2064 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04081 3115 3552 2994 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04080 2994 3114 3115 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04079 8185 3553 2994 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04078 3112 3115 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04077 2588 2733 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04076 2587 2734 2732 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04075 2586 2735 2728 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04074 8185 2964 2586 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04073 8185 3834 2735 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04072 2734 2735 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04071 8185 3267 2733 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04070 2732 2735 2588 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04069 2729 2732 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04068 8185 2729 2587 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04067 2728 2734 2729 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04066 2964 2728 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04065 8185 2728 2964 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04064 6723 6877 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04063 6722 6879 6876 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04062 6721 6878 6872 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04061 8185 6870 6721 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04060 8185 8166 6878 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04059 6879 6878 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04058 8185 6882 6877 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04057 6876 6878 6723 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04056 6873 6876 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04055 8185 6873 6722 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04054 6872 6879 6873 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04053 6870 6872 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04052 8185 6872 6870 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04051 1790 1890 1662 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04050 1662 1795 1790 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04049 8185 3150 1662 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04048 6071 6801 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04047 8185 6349 6071 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04046 6071 6549 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04045 8185 6076 6071 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04044 6070 6520 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04043 8185 6292 6070 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04042 6070 6792 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04041 8185 6541 6070 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04040 410 1115 515 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04039 515 1114 411 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04038 411 514 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04037 409 512 515 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04036 8185 1110 409 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04035 8185 517 410 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04034 1761 515 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04033 8185 3819 3614 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04032 3614 6143 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04031 3613 3614 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04030 4726 4725 4729 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04029 4729 4728 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04028 4727 6341 4726 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04027 4745 7352 4743 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04026 4743 5467 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04025 4744 4742 4745 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04024 6254 8179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04023 6415 7302 6254 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04022 8185 6418 6415 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04021 4136 4134 4135 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04020 4135 5633 4136 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04019 8185 4418 4135 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04018 4133 4136 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04017 6284 5003 4229 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04016 4229 4228 6284 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04015 8185 5908 4229 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_04014 8185 4644 3274 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04013 3274 3275 3273 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04012 3751 3273 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_04011 1230 1343 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04010 1229 1344 1342 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04009 1228 1345 1338 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04008 8185 5443 1228 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04007 8185 1772 1345 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04006 1344 1345 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_04005 8185 1526 1343 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_04004 1342 1345 1230 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04003 1339 1342 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04002 8185 1339 1229 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04001 1338 1344 1339 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_04000 5443 1338 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03999 8185 1338 5443 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03998 650 652 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03997 630 651 648 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03996 629 653 647 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03995 8185 6520 629 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03994 8185 3708 653 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03993 651 653 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03992 8185 654 652 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03991 648 653 650 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03990 649 648 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03989 8185 649 630 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03988 647 651 649 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03987 6520 647 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03986 8185 647 6520 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03985 4787 4795 4789 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03984 4789 6417 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03983 4788 4786 4787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03982 1095 1123 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03981 1332 5641 1095 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03980 1149 1148 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03979 2695 3608 1149 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03978 2905 3378 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03977 2904 3373 2905 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03976 1057 1060 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03975 1059 1061 1058 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03974 1054 1062 1055 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03973 8185 5394 1054 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03972 8185 1951 1062 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03971 1061 1062 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03970 8185 1307 1060 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03969 1058 1062 1057 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03968 1056 1058 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03967 8185 1056 1059 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03966 1055 1061 1056 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03965 5394 1055 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03964 8185 1055 5394 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03963 8185 7343 7180 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03962 7180 7342 7341 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03961 7334 7341 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03960 8185 6540 6537 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03959 6537 6536 6538 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03958 6535 6538 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03957 2089 6359 2088 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03956 2088 2217 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03955 2216 2924 2089 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03954 2090 4574 2091 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03953 2091 4302 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03952 2217 2690 2090 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03951 1554 4540 1555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03950 1555 1553 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03949 1889 1559 1554 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03948 833 4302 834 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03947 834 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03946 1361 2262 833 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03945 8185 6102 6106 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03944 6108 6823 6101 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03943 6105 7352 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_03942 6101 6100 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03941 8185 6102 6100 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_03940 6829 6108 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_03939 6106 6103 6104 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03938 6104 7352 6108 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03937 6108 6105 6107 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03936 6107 7528 6106 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03935 7687 7880 7688 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03934 7688 8179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03933 8172 7882 7687 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03932 7693 8187 7694 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03931 7694 7888 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03930 7889 8184 7693 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03929 2566 2894 2565 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03928 2565 2703 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03927 2722 4306 2566 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03926 2549 4574 2550 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03925 2550 4573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03924 3150 6293 2549 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03923 4472 4583 4378 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03922 4378 5038 4472 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03921 8185 4582 4378 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03920 8185 4424 3455 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03919 3455 3763 3573 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03918 3571 3573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03917 6551 6797 6552 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03916 6552 6802 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03915 6550 7353 6551 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03914 7541 6549 6550 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03913 8185 1133 1134 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03912 8185 1145 1134 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03911 1134 5176 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03910 1132 1134 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03909 7054 7354 7055 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03908 7055 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03907 7052 7051 7054 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03906 7053 8086 7052 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03905 4875 6636 4874 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03904 4874 6652 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03903 4873 6421 4875 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03902 5038 6921 4873 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03901 4304 4575 4305 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03900 4305 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03899 4303 6609 4304 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03898 4579 4302 4303 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03897 4872 6396 4871 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03896 4871 6636 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03895 4870 6421 4872 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03894 5037 6921 4870 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03893 3761 4172 3760 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03892 3760 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03891 3759 8139 3761 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03890 7455 7749 7457 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03889 7457 7518 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03888 7456 7725 7455 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03887 7730 7496 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03886 7496 7724 7456 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03885 8185 6396 4857 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03884 4857 7633 5014 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03883 5013 5014 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03882 7049 7354 7050 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03881 7050 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03880 7047 7353 7049 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03879 7048 8071 7047 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03878 1586 4518 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03877 8185 2698 1586 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03876 1586 5148 1587 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03875 1587 2926 1586 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03874 8185 1892 2025 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03873 8185 2700 2025 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03872 2025 1893 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03871 2942 2025 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03870 2844 3759 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03869 2843 4166 2844 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03868 8185 4510 2843 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03867 3722 3720 3721 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03866 3721 4492 3722 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03865 8185 8064 3721 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03864 6057 6489 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03863 6056 6480 6057 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03862 8185 6055 6056 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03861 6786 6056 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03860 3358 4556 3357 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03859 3357 3610 3358 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03858 8185 3788 3357 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03857 3356 3358 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03856 8185 786 785 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03855 4068 785 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03854 8185 785 4068 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03853 8185 785 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03852 8144 785 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03851 8185 786 787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03850 4573 787 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03849 8185 787 4573 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03848 8185 787 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03847 8144 787 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03846 8185 576 577 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03845 786 577 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03844 8185 577 786 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03843 8185 577 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03842 8144 577 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03841 8185 3179 2489 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03840 6543 2489 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03839 8185 2489 6543 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03838 8185 2489 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03837 8144 2489 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03836 8185 3179 2726 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03835 6797 2726 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03834 8185 2726 6797 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03833 8185 2726 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03832 8144 2726 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03831 8185 3179 2720 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03830 7356 2720 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03829 8185 2720 7356 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03828 8185 2720 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03827 8144 2720 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03826 8185 3179 3180 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03825 4051 3180 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03824 8185 3180 4051 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03823 8185 3180 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03822 8144 3180 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03821 8185 2490 2491 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03820 3179 2491 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03819 8185 2491 3179 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03818 8185 2491 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03817 8144 2491 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03816 8185 1150 430 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03815 430 3622 552 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03814 551 552 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03813 8185 1317 1218 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03812 1218 5641 1318 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03811 1956 1318 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03810 6250 6921 6251 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03809 6251 6658 6411 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03808 8185 7130 6250 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03807 6410 6411 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03806 8185 7051 2572 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03805 2572 2719 2716 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03804 2938 2716 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03803 6518 7073 6519 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03802 6519 6835 6518 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03801 8185 6794 6519 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03800 6517 6518 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03799 5338 5483 5340 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03798 5340 5654 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03797 5339 7353 5338 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03796 7880 5484 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03795 5484 7500 5339 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03794 8185 4311 3417 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03793 3417 3415 3420 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03792 3416 3420 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03791 2447 6543 2450 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03790 2450 6802 2449 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03789 8185 2687 2447 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03788 2696 2449 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03787 4209 4212 4211 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03786 4211 4208 4210 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03785 8185 4206 4209 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03784 4207 4210 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03783 6129 6131 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03782 6023 6025 6024 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03781 6021 6130 6125 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03780 8185 6127 6021 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03779 8185 7821 6130 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03778 6025 6130 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03777 8185 6128 6131 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03776 6024 6130 6129 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03775 6022 6024 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03774 8185 6022 6023 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03773 6125 6025 6022 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03772 6127 6125 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03771 8185 6125 6127 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03770 1164 5624 1165 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03769 1165 1565 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03768 1163 5483 1164 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03767 1381 1162 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03766 1162 3857 1163 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03765 2687 1799 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03764 2690 5940 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03763 774 2964 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03762 7581 7845 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03761 7270 7572 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03760 7076 7272 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03759 7617 8186 7616 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03758 7616 7619 7618 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03757 8185 7869 7617 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03756 7887 7618 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03755 3235 5147 3237 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03754 3237 4228 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03753 3236 7343 3235 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03752 3794 3346 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03751 3346 5148 3236 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03750 3922 7026 3923 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03749 3923 4573 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03748 3921 4572 3922 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03747 6090 4027 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03746 4027 5003 3921 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03745 3893 4143 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03744 4155 3986 3893 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03743 807 882 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03742 806 883 880 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03741 805 884 877 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03740 8185 1304 805 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03739 8185 1951 884 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03738 883 884 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03737 8185 885 882 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03736 880 884 807 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03735 879 880 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03734 8185 879 806 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03733 877 883 879 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03732 1304 877 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03731 8185 877 1304 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03730 7370 7779 7195 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03729 7195 7778 7370 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03728 8185 7863 7195 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03727 7367 7370 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03726 5653 6883 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03725 4134 5563 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03724 2789 5387 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03723 5380 5394 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03722 369 1799 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03721 8185 2492 369 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03720 579 2968 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03719 8185 2964 579 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03718 1901 2471 1903 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03717 1903 1902 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03716 1900 1899 1901 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03715 3642 2033 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03714 2033 2035 1900 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03713 3230 3316 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03712 3546 3229 3230 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03711 8164 8168 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03710 8163 8167 8165 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03709 8160 8170 8161 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03708 8185 8159 8160 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03707 8185 8166 8170 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03706 8167 8170 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03705 8185 8173 8168 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03704 8165 8170 8164 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03703 8162 8165 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03702 8185 8162 8163 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03701 8161 8167 8162 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03700 8159 8161 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03699 8185 8161 8159 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03698 7044 7041 7042 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03697 7042 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03696 7043 8071 7044 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03695 5156 7056 5157 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03694 5157 6294 5156 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03693 8185 5162 5157 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03692 5416 5156 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03691 8185 2906 2004 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03690 2004 2011 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03689 2005 2004 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03688 8185 2906 2002 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03687 2002 2006 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03686 2003 2002 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03685 1227 5641 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03684 1346 1335 1227 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03683 7729 7955 7168 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03682 7168 7747 7729 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03681 8185 7319 7168 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03680 3234 3763 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03679 3327 4424 3234 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03678 6682 6773 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03677 6681 6774 6772 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03676 6680 6776 6768 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03675 8185 6775 6680 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03674 8185 8063 6776 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03673 6774 6776 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03672 8185 6780 6773 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03671 6772 6776 6682 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03670 6770 6772 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03669 8185 6770 6681 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03668 6768 6774 6770 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03667 6775 6768 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03666 8185 6768 6775 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03665 6093 6095 6094 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03664 8185 6094 6319 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03663 8185 6095 6097 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03662 6092 6096 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03661 6094 6097 6092 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03660 8185 6344 6093 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03659 6319 6094 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03658 5765 5842 5918 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03657 8185 5918 6096 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03656 8185 5842 5844 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03655 5766 7549 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03654 5918 5844 5766 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03653 8185 6292 5765 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03652 6096 5918 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03651 5132 7787 5127 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03650 5127 5907 5132 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03649 8185 6076 5127 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03648 1575 2469 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03647 2924 7051 1575 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03646 1211 5828 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03645 1306 1313 1211 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03644 2212 2894 2086 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03643 2085 7051 2212 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03642 2086 4067 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03641 2679 2212 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03640 8185 2210 2085 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03639 2085 2682 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03638 2389 4947 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03637 2648 3134 2389 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03636 8131 8133 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03635 8129 8134 8132 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03634 8126 8135 8127 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03633 8185 8125 8126 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03632 8185 8166 8135 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03631 8134 8135 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03630 8185 8130 8133 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03629 8132 8135 8131 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03628 8128 8132 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03627 8185 8128 8129 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03626 8127 8134 8128 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03625 8125 8127 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03624 8185 8127 8125 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03623 8185 6785 6059 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03622 6059 6784 6058 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03621 6503 6058 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03620 8185 5616 5297 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03619 5297 5414 5407 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03618 6785 5407 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03617 8185 7352 6547 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03616 6547 7883 6548 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03615 7760 6548 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03614 6122 6362 6356 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03613 8185 6356 6581 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03612 8185 6362 6357 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03611 6126 6576 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03610 6356 6357 6126 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03609 8185 6353 6122 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03608 6581 6356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03607 6117 6359 6119 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03606 8185 6119 6353 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03605 8185 6359 6120 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03604 6121 7777 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03603 6119 6120 6121 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03602 8185 6347 6117 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_03601 6353 6119 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03600 1261 2469 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03599 1996 4306 1261 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03598 7637 7888 7638 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03597 7638 7643 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03596 7877 7891 7637 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03595 7018 7352 7019 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03594 7019 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03593 7017 8021 7018 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03592 2799 3581 2800 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03591 2800 3586 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03590 2797 2796 2799 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03589 2798 3542 2797 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03588 3003 3146 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03587 3143 4007 3003 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03586 8185 4510 3143 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03585 1916 1918 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03584 1879 1917 1878 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03583 1876 1919 1913 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03582 8185 5906 1876 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03581 8185 3708 1919 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03580 1917 1919 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03579 8185 3508 1918 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03578 1878 1919 1916 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03577 1877 1878 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03576 8185 1877 1879 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03575 1913 1917 1877 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03574 5906 1913 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03573 8185 1913 5906 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03572 7312 7518 7162 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03571 7162 7313 7312 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03570 8185 7314 7162 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03569 7486 7312 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03568 4653 6792 4652 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03567 4652 5384 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03566 4651 5606 4653 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03565 5551 5888 5550 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03564 8185 7500 5552 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03563 5550 5552 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03562 3395 5483 3394 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03561 3394 5654 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03560 3396 6293 3395 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03559 3393 4461 3396 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03558 2516 4172 2517 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03557 2517 4173 2615 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03556 8185 7585 2516 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03555 2614 2615 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03554 8185 4022 4023 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03553 6152 4023 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03552 8185 4023 6152 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03551 8185 4023 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03550 8144 4023 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03549 8185 3792 3793 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03548 5961 3793 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03547 8185 3793 5961 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03546 8185 3793 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03545 8144 3793 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03544 8185 6152 6153 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03543 8166 6153 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03542 8185 6153 8166 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03541 8185 6153 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03540 8144 6153 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03539 8185 6152 6151 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03538 7821 6151 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03537 8185 6151 7821 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03536 8185 6151 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03535 8144 6151 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03534 8185 6152 5963 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03533 5864 5963 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03532 8185 5963 5864 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03531 8185 5963 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03530 8144 5963 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03529 8185 5961 5962 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03528 5863 5962 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03527 8185 5962 5863 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03526 8185 5962 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03525 8144 5962 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03524 8185 6152 6069 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03523 8063 6069 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03522 8185 6069 8063 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03521 8185 6069 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03520 8144 6069 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03519 8185 6152 6068 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03518 6067 6068 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03517 8185 6068 6067 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03516 8185 6068 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03515 8144 6068 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03514 1445 1447 5558 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03513 8185 5453 1445 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03512 1444 1446 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03511 5558 1443 1444 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03510 8185 1446 1447 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03509 1443 5453 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03508 8185 8175 8177 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03507 8177 8182 8178 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03506 8176 8178 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03505 8185 4955 4232 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03504 4231 4232 4233 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03503 8185 4230 4231 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03502 4530 4233 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03501 8185 4233 4530 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03500 8185 2968 792 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03499 790 792 789 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03498 8185 2964 790 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03497 791 789 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03496 8185 789 791 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03495 2960 2958 2959 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03494 2959 3860 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03493 3073 2957 2960 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03492 3484 5483 3483 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03491 3483 5654 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03490 3482 6293 3484 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03489 3622 5015 3482 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03488 2515 3566 2514 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03487 2514 3293 2613 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03486 8185 3744 2515 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03485 2612 2613 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03484 3732 4167 3733 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03483 3733 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03482 3731 6796 3732 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03481 3730 6273 3731 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03480 5909 5603 5604 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03479 8185 7314 5605 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03478 5604 5605 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03477 5709 6632 5708 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03476 5708 7633 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03475 5707 5868 5709 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03474 5706 7130 5707 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03473 6617 6629 6616 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03472 6616 6615 6617 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03471 8185 6614 6616 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03470 8185 4647 4650 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03469 4650 5379 4649 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03468 4648 4649 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03467 4938 5429 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03466 8185 7787 4938 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03465 4938 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03464 8185 8045 4938 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03463 4934 4938 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03462 3480 3621 3639 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03461 8185 5453 3480 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03460 3481 3787 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03459 3639 3619 3481 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03458 8185 3787 3621 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03457 3619 5453 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03456 4825 4922 4924 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03455 8185 7056 4825 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03454 4826 4921 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03453 4924 4919 4826 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03452 8185 4921 4922 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03451 4919 7056 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03450 7552 7804 7551 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03449 7553 7550 7552 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03448 7551 7554 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03447 7547 7552 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03446 8185 7548 7553 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03445 7553 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_03444 8185 5408 5137 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03443 5137 5140 5138 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03442 5136 5138 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03441 8185 5168 3471 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03440 3471 3608 3609 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03439 3801 3609 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03438 8185 5147 1658 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03437 1658 4228 1781 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03436 1780 1781 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03435 8185 2968 442 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03434 442 2964 575 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03433 574 575 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03432 8185 2718 2458 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03431 2458 2719 2459 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03430 2706 2459 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03429 6066 8008 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03428 6301 6285 6066 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03427 6065 6286 6301 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03426 8185 6267 6065 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03425 6064 6520 6301 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03424 8185 6284 6064 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03423 3306 3987 3305 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03422 3305 3993 3306 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03421 8185 3315 3305 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03420 3303 3306 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03419 4005 7056 3908 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03418 3908 5406 4005 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03417 8185 6812 3908 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03416 4003 4005 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03415 2409 2413 2410 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03414 2410 2886 2411 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03413 8185 2407 2409 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03412 2408 2411 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03411 6713 6846 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03410 6712 6848 6845 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03409 6711 6847 6840 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03408 8185 6838 6711 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03407 8185 7821 6847 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03406 6848 6847 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03405 8185 6843 6846 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03404 6845 6847 6713 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03403 6841 6845 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03402 8185 6841 6712 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03401 6840 6848 6841 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03400 6838 6840 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03399 8185 6840 6838 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03398 6727 6890 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03397 6726 6892 6889 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03396 6725 6891 6885 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03395 8185 6883 6725 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03394 8185 8166 6891 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03393 6892 6891 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03392 8185 6899 6890 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03391 6889 6891 6727 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03390 6886 6889 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03389 8185 6886 6726 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03388 6885 6892 6886 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03387 6883 6885 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03386 8185 6885 6883 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03385 4721 4722 4723 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03384 4723 7352 4721 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03383 8185 4739 4723 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03382 5344 6900 5345 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03381 5345 8187 5493 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03380 8185 7883 5344 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03379 5492 5493 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03378 7407 7881 7221 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03377 7221 7408 7407 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03376 8185 7891 7221 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03375 7305 7407 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03374 3000 3582 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03373 3133 3356 3000 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03372 8185 3579 3133 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03371 3552 3133 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03370 2171 4189 2062 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03369 2062 2170 2171 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03368 8185 2375 2062 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03367 2168 2171 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03366 667 669 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03365 633 668 665 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03364 632 670 664 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03363 8185 677 632 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03362 8185 1951 670 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03361 668 670 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03360 8185 671 669 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03359 665 670 667 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03358 666 665 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03357 8185 666 633 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03356 664 668 666 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03355 677 664 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03354 8185 664 677 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03353 8185 7774 8006 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03352 8006 7767 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03351 8185 7768 8006 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03350 1052 1743 1053 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03349 1053 1744 1052 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03348 8185 8045 1053 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03347 1606 4295 1607 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03346 1607 4310 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03345 1604 4293 1606 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03344 1897 1605 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_03343 1605 5648 1604 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03342 4640 5737 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03341 4802 5740 4640 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03340 7649 7738 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03339 7728 7730 7649 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03338 2318 5453 1192 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03337 8185 7314 1282 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03336 1192 1282 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03335 6236 6393 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03334 6235 6395 6390 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03333 6234 6394 6388 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03332 8185 6398 6234 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03331 8185 8166 6394 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03330 6395 6394 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03329 8185 6401 6393 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03328 6390 6394 6236 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03327 6391 6390 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03326 8185 6391 6235 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03325 6388 6395 6391 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03324 6398 6388 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03323 8185 6388 6398 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03322 6665 7884 6666 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03321 6666 7408 6665 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03320 8185 7891 6666 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03319 6914 6665 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03318 2172 2179 1960 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03317 1960 2178 2172 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03316 8185 3148 1960 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03315 2388 3780 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03314 3556 4255 2388 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03313 2829 3990 2828 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03312 2828 3989 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03311 2827 3348 2829 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03310 2071 2190 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03309 2072 2191 2188 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03308 2070 2192 2184 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03307 8185 5143 2070 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03306 8185 3708 2192 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03305 2191 2192 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03304 8185 2189 2190 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03303 2188 2192 2071 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03302 2185 2188 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03301 8185 2185 2072 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03300 2184 2191 2185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03299 5143 2184 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03298 8185 2184 5143 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03297 640 1123 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03296 903 1115 640 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03295 3254 3624 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03294 3629 3253 3254 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03293 7656 7754 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03292 7743 7742 7656 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03291 3896 4172 3897 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03290 3897 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03289 3989 7349 3896 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03288 2982 3088 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03287 2981 3083 3085 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03286 2980 3091 3081 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03285 8185 6792 2980 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03284 8185 3708 3091 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03283 3083 3091 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03282 8185 3962 3088 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03281 3085 3091 2982 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03280 3084 3085 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03279 8185 3084 2981 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03278 3081 3083 3084 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03277 6792 3081 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03276 8185 3081 6792 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03275 8185 7343 6213 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03274 6213 6298 6299 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03273 6297 6299 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03272 5360 6909 5359 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03271 5359 5971 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03270 5502 7633 5360 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03269 641 1123 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03268 939 1114 641 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03267 2559 4068 2560 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03266 2560 6311 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03265 2693 6293 2559 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03264 5239 6652 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03263 5238 6172 5239 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03262 8185 3556 1645 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03261 1735 2672 1642 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03260 1733 3958 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_03259 1642 1730 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03258 8185 3556 1730 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_03257 1729 1735 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_03256 1645 1732 1643 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03255 1643 3958 1735 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03254 1735 1733 1644 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03253 1644 2155 1645 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03252 8185 3556 1939 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03251 1941 3009 1934 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03250 1938 3958 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_03249 1934 1935 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03248 8185 3556 1935 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_03247 2132 1941 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_03246 1939 1936 1937 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03245 1937 3958 1941 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03244 1941 1938 1940 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03243 1940 2154 1939 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03242 8185 3990 2991 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03241 2991 3989 3105 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03240 3104 3105 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03239 1516 1515 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03238 1513 1517 1514 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03237 1511 1518 1510 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03236 8185 5419 1511 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03235 8185 1772 1518 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03234 1517 1518 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_03233 8185 1519 1515 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_03232 1514 1518 1516 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03231 1512 1514 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03230 8185 1512 1513 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03229 1510 1517 1512 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03228 5419 1510 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03227 8185 1510 5419 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03226 5081 6478 5083 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03225 5083 6477 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03224 5082 6472 5081 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03223 7318 6473 5082 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03222 3076 6472 2978 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03221 2978 6473 3076 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03220 8185 8064 2978 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03219 6087 3076 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03218 5726 6921 5725 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03217 5725 6176 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03216 5724 7130 5726 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03215 7264 7835 7233 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03214 8185 7957 7265 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03213 7233 7265 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03212 3414 4575 3413 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03211 3413 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03210 3412 6609 3414 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03209 4582 4306 3412 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03208 6652 7398 6653 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03207 6653 7884 6652 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03206 8185 7891 6653 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03205 1752 1965 1219 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03204 1219 1964 1752 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03203 8185 3148 1219 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03202 2015 4172 2016 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03201 2016 4173 2014 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03200 8185 7549 2015 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03199 2156 2014 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03198 8185 3556 1636 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03197 1715 3958 1633 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03196 1714 2144 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_03195 1633 1712 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03194 8185 3556 1712 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_03193 1711 1715 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_03192 1636 1925 1634 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03191 1634 2144 1715 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03190 1715 1714 1635 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03189 1635 2605 1636 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03188 8185 3556 1464 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03187 1463 1467 1458 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03186 1461 2144 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_03185 1458 1459 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03184 8185 3556 1459 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_03183 2136 1463 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_03182 1464 1932 1460 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03181 1460 2144 1463 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03180 1463 1461 1462 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03179 1462 2608 1464 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_03178 7189 7354 7190 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03177 7190 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03176 7188 7353 7189 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03175 7342 7824 7188 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03174 2927 2926 2928 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03173 2928 2924 2927 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03172 8185 2925 2928 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03171 3405 2927 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03170 7004 7002 7003 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03169 7003 7250 7005 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03168 8185 7011 7004 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03167 7508 7005 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03166 1682 1891 1681 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03165 1681 1796 1797 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03164 8185 6363 1682 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03163 4236 1797 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03162 8185 1806 1666 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03161 1666 2926 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03160 2232 1805 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03159 1666 2924 1805 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03158 1805 2698 1666 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03157 8185 3251 3392 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03156 8185 3250 3392 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03155 3392 3252 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03154 3409 3392 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03153 5838 6090 5763 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03152 5763 6089 5838 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03151 8185 6344 5763 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03150 2985 3093 3720 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03149 8185 3095 2985 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03148 2986 3100 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03147 3720 3094 2986 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03146 8185 3100 3093 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03145 3094 3095 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03144 8185 4076 3855 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03143 7026 3855 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03142 8185 3855 7026 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03141 8185 3855 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03140 8144 3855 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03139 8185 4076 4077 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03138 6609 4077 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03137 8185 4077 6609 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03136 8185 4077 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03135 8144 4077 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03134 8185 4076 4065 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03133 7354 4065 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03132 8185 4065 7354 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03131 8185 4065 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03130 8144 4065 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03129 8185 3662 3663 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03128 4076 3663 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03127 8185 3663 4076 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03126 8185 3663 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03125 8144 3663 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03124 8185 568 567 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03123 4293 567 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03122 8185 567 4293 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03121 8185 567 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03120 8144 567 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03119 8185 568 569 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03118 4302 569 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03117 8185 569 4302 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03116 8185 569 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03115 8144 569 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03114 8185 568 566 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03113 4572 566 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03112 8185 566 4572 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03111 8185 566 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03110 8144 566 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03109 8185 375 376 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03108 568 376 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03107 8185 376 568 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03106 8185 376 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03105 8144 376 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03104 5922 5653 5643 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03103 5643 5641 5922 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03102 8185 5642 5643 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03101 8185 5728 5715 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03100 5715 5870 5716 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03099 5967 5716 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03098 6742 7884 6741 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03097 6741 7398 6910 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03096 8185 7883 6742 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03095 6909 6910 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03094 7532 7750 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03093 8185 7787 7532 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03092 7532 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03091 8185 8045 7532 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03090 7566 7532 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03089 4515 6304 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03088 8185 7787 4515 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03087 4515 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03086 8185 8045 4515 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_03085 4433 4515 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03084 7736 7734 7653 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03083 7653 7962 7736 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03082 8185 7957 7653 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03081 7733 7736 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03080 8185 782 571 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03079 4306 571 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03078 8185 571 4306 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03077 8185 571 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03076 8144 571 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03075 8185 782 570 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03074 4067 570 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03073 8185 570 4067 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03072 8185 570 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03071 8144 570 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03070 8185 782 783 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03069 5624 783 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03068 8185 783 5624 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03067 8185 783 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03066 8144 783 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03065 8185 378 377 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03064 782 377 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03063 8185 377 782 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03062 8185 377 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03061 8144 377 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03060 8185 1190 1191 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03059 4574 1191 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03058 8185 1191 4574 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03057 8185 1191 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03056 8144 1191 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03055 8185 1190 971 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03054 5648 971 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03053 8185 971 5648 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03052 8185 971 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03051 8144 971 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03050 8185 1190 967 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03049 4167 967 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03048 8185 967 4167 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03047 8185 967 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03046 8144 967 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03045 8185 791 788 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03044 1190 788 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03043 8185 788 1190 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03042 8185 788 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03041 8144 788 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03040 6477 6304 6215 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03039 6215 7747 6477 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03038 8185 6535 6215 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03037 6635 7408 6637 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03036 6637 7892 6638 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03035 8185 7883 6635 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03034 6654 6638 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_03033 8185 2233 2100 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03032 2100 2232 2231 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03031 2240 2231 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03030 8185 4306 2470 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03029 2470 2469 2472 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03028 2943 2472 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03027 8185 2723 2582 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03026 2582 2722 2724 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03025 3415 2724 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03024 8185 4049 3825 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03023 4295 3825 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03022 8185 3825 4295 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03021 8185 3825 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03020 8144 3825 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03019 8185 4049 4050 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03018 4575 4050 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03017 8185 4050 4575 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03016 8185 4050 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03015 8144 4050 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03014 8185 4045 4046 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03013 4049 4046 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03012 8185 4046 4049 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03011 8185 4046 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03010 8144 4046 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03009 7369 7059 7060 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03008 7060 7058 7369 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03007 8185 7062 7060 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_03006 8185 2227 2018 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03005 2018 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03004 2235 2017 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03003 2018 2203 2017 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03002 2017 2926 2018 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_03001 8185 8184 5789 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_03000 5789 7893 5974 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02999 5878 5974 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02998 8185 4574 2443 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02997 2443 4068 2444 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02996 2688 2444 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02995 1272 4067 1273 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02994 1273 2719 1386 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02993 8185 3857 1272 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02992 1389 1386 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02991 346 1150 345 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02990 345 359 347 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02989 8185 4558 346 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02988 343 347 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02987 7960 7954 6467 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02986 8185 8064 6468 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02985 6467 6468 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02984 1082 1086 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02983 1084 1085 1083 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02982 1079 1087 1080 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02981 8185 1758 1079 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02980 8185 1772 1087 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02979 1085 1087 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02978 8185 1091 1086 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02977 1083 1087 1082 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02976 1081 1083 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02975 8185 1081 1084 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02974 1080 1085 1081 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02973 1758 1080 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02972 8185 1080 1758 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02971 8185 6618 5682 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02970 5682 6398 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02969 8185 6141 5682 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02968 8185 6127 5665 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02967 5665 5664 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02966 8185 6143 5665 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02965 4541 4987 4353 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02964 4353 4749 4541 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02963 8185 4540 4353 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02962 4449 4541 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02961 6736 7619 6737 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02960 6737 6907 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02959 6735 8186 6736 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02958 6906 6908 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02957 6908 8184 6735 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02956 5634 5632 5635 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02955 5635 5633 5634 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02954 8185 7547 5635 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02953 5912 5634 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02952 5129 5419 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02951 5567 5571 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02950 5632 5435 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02949 2608 2809 2512 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02948 2512 3320 2608 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02947 8185 3315 2512 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02946 2831 2833 2832 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02945 2832 3310 2831 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02944 8185 2830 2832 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02943 4498 2831 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02942 5782 5957 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02941 5781 5958 5955 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02940 5780 5960 5952 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02939 8185 6143 5780 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02938 8185 7821 5960 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02937 5958 5960 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02936 8185 6386 5957 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02935 5955 5960 5782 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02934 5954 5955 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02933 8185 5954 5781 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02932 5952 5958 5954 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02931 6143 5952 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02930 8185 5952 6143 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02929 8185 2439 1795 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02928 1795 1792 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02927 8185 2003 1795 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02926 817 3608 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02925 948 1372 817 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02924 5444 5443 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02923 5421 5143 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02922 7758 7979 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02921 8009 8008 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02920 7955 7954 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02919 7802 3077 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02918 1277 4293 1278 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02917 1278 4068 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02916 1276 4574 1277 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02915 1617 1393 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02914 1393 4075 1276 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02913 2114 6797 2115 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02912 2115 4575 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02911 2113 4306 2114 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02910 2254 2255 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02909 2255 5942 2113 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02908 3749 4511 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02907 3748 4512 3749 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02906 1103 1102 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02905 1100 1104 1101 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02904 1098 1105 1097 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02903 8185 1335 1098 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02902 8185 1772 1105 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02901 1104 1105 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02900 8185 1330 1102 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02899 1101 1105 1103 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02898 1099 1101 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02897 8185 1099 1100 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02896 1097 1104 1099 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02895 1335 1097 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02894 8185 1097 1335 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02893 4365 4566 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02892 4366 4567 4565 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02891 4364 4569 4564 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02890 8185 4734 4364 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02889 8185 5864 4569 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02888 4567 4569 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02887 8185 4570 4566 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02886 4565 4569 4365 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02885 4568 4565 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02884 8185 4568 4366 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02883 4564 4567 4568 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02882 4734 4564 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02881 8185 4564 4734 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02880 3372 4302 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02879 8185 5624 3372 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02878 3372 3370 4529 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02877 4529 3371 3372 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02876 4396 4537 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02875 4963 4727 4396 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02874 4636 6383 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02873 4766 4635 4636 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02872 4730 4230 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02871 4193 4021 3773 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02870 3773 7788 4193 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02869 8185 6792 3773 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02868 1914 6867 2129 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02867 8185 2129 2126 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02866 8185 6867 2131 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02865 1915 2133 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02864 2129 2131 1915 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02863 8185 2127 1914 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02862 2126 2129 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02861 2362 4685 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02860 3562 2361 2362 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02859 7185 7352 7184 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02858 7184 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02857 7336 7824 7185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02856 6116 6358 6352 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02855 8185 6352 6347 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02854 8185 6358 6350 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02853 6118 6349 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02852 6352 6350 6118 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02851 8185 6586 6116 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02850 6347 6352 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02849 2936 5496 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02848 2935 4790 2936 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02847 1675 4437 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02846 1753 1752 1675 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02845 2528 2635 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02844 2636 3137 2528 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02843 1289 1451 1196 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02842 1195 1929 1289 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02841 1196 2132 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02840 1296 1289 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02839 8185 1287 1195 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02838 1195 2595 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02837 6496 6497 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02836 6493 6498 6494 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02835 6491 6499 6490 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02834 8185 6489 6491 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02833 8185 8063 6499 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02832 6498 6499 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02831 8185 6495 6497 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02830 6494 6499 6496 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02829 6492 6494 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02828 8185 6492 6493 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02827 6490 6498 6492 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02826 6489 6490 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02825 8185 6490 6489 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02824 4537 4234 4235 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02823 4235 4447 4537 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02822 8185 5449 4235 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02821 6146 6383 6376 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02820 8185 6376 6374 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02819 8185 6383 6379 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02818 6147 6378 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02817 6376 6379 6147 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02816 8185 6375 6146 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02815 6374 6376 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02814 4810 7887 4811 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02813 4811 6421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02812 5042 7149 4810 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02811 4829 5600 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02810 4929 4927 4829 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02809 1881 4228 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02808 2199 5147 1881 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02807 3791 7354 3790 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02806 3790 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02805 3789 7353 3791 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02804 3788 3787 3789 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02803 8112 8115 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02802 8114 8116 8113 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02801 8108 8117 8110 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02800 8185 8119 8108 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02799 8185 8166 8117 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02798 8116 8117 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02797 8185 8118 8115 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02796 8113 8117 8112 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02795 8111 8113 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02794 8185 8111 8114 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02793 8110 8116 8111 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02792 8119 8110 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02791 8185 8110 8119 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02790 8185 7796 7665 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02789 7665 7794 7795 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02788 7793 7795 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02787 5589 5588 5590 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02786 5590 6785 5589 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02785 8185 5587 5590 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02784 5657 5654 5656 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02783 5656 5854 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02782 5655 5942 5657 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02781 5927 6796 5655 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02780 5336 7871 5481 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02779 8185 5481 5478 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02778 8185 7871 5482 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02777 5337 5712 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02776 5481 5482 5337 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02775 8185 5664 5336 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02774 5478 5481 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02773 4256 7871 4258 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02772 8185 4258 4254 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02771 8185 7871 4259 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02770 4257 5013 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02769 4258 4259 4257 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02768 8185 4255 4256 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02767 4254 4258 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02766 4763 7871 4762 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02765 8185 4762 4759 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02764 8185 7871 4764 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02763 4761 5495 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02762 4762 4764 4761 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02761 8185 4760 4763 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02760 4759 4762 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02759 8185 7137 5723 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02758 5721 5723 5722 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02757 8185 5968 5721 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02756 5720 5722 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02755 8185 5722 5720 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02754 3333 3581 3335 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02753 3335 3356 3334 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02752 8185 3582 3333 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02751 3744 3334 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02750 5198 7871 5199 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02749 8185 5199 5196 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02748 8185 7871 5200 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02747 5201 6154 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02746 5199 5200 5201 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02745 8185 5197 5198 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02744 5196 5199 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02743 7782 7020 7021 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02742 7021 7058 7782 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02741 8185 7025 7021 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02740 8185 1381 1382 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02739 1382 1384 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02738 2249 1382 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02737 8185 1168 1166 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02736 1166 1169 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02735 1589 1166 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02734 3171 1571 1572 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02733 1572 1570 3171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02732 8185 7550 1572 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02731 7138 7888 7139 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02730 7139 7884 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02729 7136 7630 7138 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02728 7137 8184 7136 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02727 4383 4790 4384 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02726 4384 5737 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02725 4476 5740 4383 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02724 756 6609 755 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02723 755 4573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02722 4228 4302 756 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02721 2013 2220 2012 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02720 2012 2011 2013 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02719 8185 8159 2012 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02718 6278 6786 6054 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02717 6054 6503 6278 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02716 8185 7500 6054 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02715 6225 6363 6362 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02714 8185 6363 6364 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02713 6226 6607 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02712 6362 6364 6226 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02711 8185 6359 6225 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02710 6013 6500 6014 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02709 6014 6051 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02708 6012 6786 6013 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02707 6473 6046 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02706 6046 6503 6012 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02705 2874 2879 2877 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02704 8185 2873 2874 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02703 2878 2875 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02702 2877 2876 2878 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02701 8185 2875 2879 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02700 2876 2873 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02699 7640 8187 7642 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02698 7642 7892 7641 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02697 8185 7891 7640 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02696 7639 7641 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02695 8185 7356 2899 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02694 2899 6802 2900 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02693 2898 2900 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02692 8185 1590 1592 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02691 1592 3253 1591 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02690 1819 1591 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02689 1143 7051 1142 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02688 1141 1140 1143 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02687 1142 2894 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02686 1139 1143 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02685 8185 1353 1141 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02684 1141 4067 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_02683 5131 5129 5130 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02682 5130 5633 5131 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02681 8185 6530 5130 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02680 5151 5131 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02679 7635 7888 7634 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02678 7634 7643 7636 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02677 8185 7891 7635 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02676 7633 7636 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02675 3058 3858 3057 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02674 3057 3260 3185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02673 8185 3184 3058 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02672 3192 3185 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02671 4029 4538 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02670 8185 4230 4029 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02669 3307 3987 3308 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02668 3308 3993 3307 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02667 8185 3315 3308 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02666 6813 7612 6704 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02665 6704 6835 6813 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02664 8185 7342 6704 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02663 6812 6813 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02662 425 545 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02661 424 546 543 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02660 423 547 540 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02659 8185 739 423 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02658 8185 3834 547 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02657 546 547 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02656 8185 740 545 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02655 543 547 425 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02654 541 543 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02653 8185 541 424 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02652 540 546 541 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02651 739 540 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02650 8185 540 739 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02649 6249 6912 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02648 6409 6407 6249 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02647 6248 7135 6409 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02646 8185 6909 6248 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02645 6247 6410 6409 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02644 8185 6647 6247 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02643 7131 7893 7133 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02642 7133 7630 7132 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02641 8185 8184 7131 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02640 7130 7132 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02639 8185 2919 3636 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02638 3636 2918 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02637 8185 3251 3636 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02636 1612 1611 1614 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02635 1614 1619 1613 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02634 8185 2448 1612 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02633 3863 1613 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02632 6717 6860 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02631 6718 6861 6859 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02630 6716 6862 6855 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02629 8185 6864 6716 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02628 8185 7821 6862 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02627 6861 6862 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02626 8185 6863 6860 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02625 6859 6862 6717 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02624 6856 6859 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02623 8185 6856 6718 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02622 6855 6861 6856 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02621 6864 6855 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02620 8185 6855 6864 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02619 4703 4704 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02618 4625 4627 4626 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02617 4623 4706 4702 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02616 8185 4714 4623 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02615 8185 8063 4706 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02614 4627 4706 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02613 8185 7549 4704 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02612 4626 4706 4703 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02611 4624 4626 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02610 8185 4624 4625 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02609 4702 4627 4624 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02608 4714 4702 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02607 8185 4702 4714 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02606 8185 7525 7772 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02605 7772 7459 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02604 8185 7529 7772 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02603 12 88 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02602 11 89 87 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02601 10 90 83 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02600 8185 268 10 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02599 8185 1951 90 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02598 89 90 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02597 8185 91 88 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02596 87 90 12 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02595 85 87 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02594 8185 85 11 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02593 83 89 85 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02592 268 83 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02591 8185 83 268 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02590 5689 5688 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02589 5686 5690 5687 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02588 5684 5691 5683 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02587 8185 6141 5684 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02586 8185 5864 5691 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02585 5690 5691 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02584 8185 5704 5688 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02583 5687 5691 5689 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02582 5685 5687 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02581 8185 5685 5686 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02580 5683 5690 5685 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02579 6141 5683 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02578 8185 5683 6141 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02577 5823 7020 5570 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02576 5570 6294 5823 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02575 8185 5825 5570 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02574 5315 5908 5316 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02573 5316 6359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02572 5923 6363 5315 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02571 8185 6145 6111 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02570 6111 6618 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02569 6112 6111 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02568 8007 8006 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02567 8015 8004 8007 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02566 6172 7881 6171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02565 6171 7408 6172 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02564 8185 7891 6171 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02563 3466 3600 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02562 3465 3601 3598 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02561 3464 3599 3593 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02560 8185 3787 3464 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02559 8185 3834 3599 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02558 3601 3599 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02557 8185 3596 3600 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02556 3598 3599 3466 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02555 3595 3598 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02554 8185 3595 3465 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02553 3593 3601 3595 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02552 3787 3593 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02551 8185 3593 3787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02550 3434 3529 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02549 3433 3531 3526 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02548 3432 3530 3523 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02547 8185 6541 3432 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02546 8185 3708 3530 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02545 3531 3530 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02544 8185 3718 3529 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02543 3526 3530 3434 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02542 3525 3526 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02541 8185 3525 3433 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02540 3523 3531 3525 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02539 6541 3523 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02538 8185 3523 6541 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02537 7727 7725 7648 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02536 7648 7724 7727 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02535 8185 7957 7648 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02534 7723 7727 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02533 6103 6112 5767 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02532 5767 5919 6103 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02531 8185 6015 5767 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02530 8173 8171 8174 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02529 8174 8172 8173 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02528 8185 8169 8174 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02527 2555 4306 2556 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02526 2556 4574 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02525 2901 2690 2555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02524 47 1150 48 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02523 48 359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02522 165 3384 47 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02521 2676 3603 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02520 8185 2887 2676 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02519 2676 2888 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02518 8185 3606 2676 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02517 2672 2676 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02516 8185 5168 2087 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02515 2087 2217 2215 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02514 2214 2215 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02513 8185 3229 2529 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02512 2529 2847 2637 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02511 2642 2637 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02510 7035 7034 7037 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02509 7037 7043 7036 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02508 8185 7038 7035 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02507 7033 7036 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02506 6079 6543 6078 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02505 6078 6311 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02504 6077 7353 6079 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02503 6307 6076 6077 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02502 6115 6358 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02501 6340 6359 6115 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02500 8185 7788 6340 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02499 8185 5178 5174 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02498 5174 5445 5175 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02497 5642 5175 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02496 6140 6161 6139 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02495 6139 6138 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02494 6137 7887 6140 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02493 1127 4293 1126 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02492 1126 6543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02491 1986 5648 1127 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02490 4639 7633 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02489 4803 7130 4639 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02488 42 553 43 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02487 43 365 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02486 344 166 42 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02485 353 1150 351 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02484 351 359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02483 352 4251 353 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02482 8185 4255 2377 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02481 2377 3780 2376 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02480 2375 2376 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02479 2508 3730 2509 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02478 2509 3735 2603 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02477 8185 3744 2508 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02476 2601 2603 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02475 6612 6609 6611 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02474 6611 7356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02473 6610 7353 6612 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02472 7062 8097 6610 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02471 832 5447 831 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02470 831 4067 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02469 1372 5942 832 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02468 1130 4228 1131 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02467 1131 3608 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02466 1129 5147 1130 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02465 1788 1128 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02464 1128 1372 1129 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02463 8185 1798 766 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02462 766 1800 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02461 763 765 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02460 766 764 765 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02459 765 7548 766 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02458 7330 7797 7175 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02457 7175 7798 7330 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02456 8185 7349 7175 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02455 8185 5154 5153 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02454 5153 5151 5152 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02453 5150 5152 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02452 8185 4934 4694 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02451 4694 5133 4695 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02450 4693 4695 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02449 2891 2890 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02448 8185 7779 2891 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02447 2891 2889 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02446 8185 7778 2891 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02445 3771 2891 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02444 8185 1905 2040 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02443 8185 1904 2040 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02442 2040 2043 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02441 2041 2040 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02440 6256 6636 6257 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02439 6257 6909 6419 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02438 8185 6921 6256 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02437 6418 6419 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02436 777 2968 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02435 8185 5940 777 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02434 777 2262 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02433 8185 2964 777 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02432 778 777 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02431 8185 2035 2038 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02430 2038 2036 2037 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02429 2485 2037 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02428 2504 2593 2794 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02427 8185 2589 2504 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02426 2505 2591 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02425 2794 2590 2505 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02424 8185 2591 2593 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02423 2590 2589 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02422 3427 5077 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02421 3510 7318 3427 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02420 8185 3507 3510 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02419 3508 3510 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02418 6163 7881 6164 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02417 6164 7398 6162 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02416 8185 8184 6163 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02415 6161 6162 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02414 8185 7130 6750 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02413 6750 6921 6919 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02412 7151 6919 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02411 8185 1372 1257 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02410 1257 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02409 1576 1370 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02408 1257 4518 1370 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02407 1370 2926 1257 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02406 5749 6273 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02405 5894 6480 5749 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02404 8185 5823 5894 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02403 6051 5894 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02402 1692 5648 1693 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02401 1693 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02400 1691 5447 1692 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02399 1905 1830 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02398 1830 7051 1691 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02397 3938 4572 3937 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02396 3937 4051 4052 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02395 8185 5483 3938 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02394 4997 4052 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02393 1071 1070 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02392 1068 1072 1067 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02391 1065 1073 1064 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02390 8185 1063 1065 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02389 8185 1951 1073 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02388 1072 1073 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02387 8185 1069 1070 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02386 1067 1073 1071 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02385 1066 1067 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02384 8185 1066 1068 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02383 1064 1072 1066 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02382 1063 1064 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02381 8185 1064 1063 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02380 5773 5934 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02379 5772 5931 5933 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02378 5771 5936 5930 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02377 8185 5938 5771 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02376 8185 7821 5936 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02375 5931 5936 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02374 8185 5935 5934 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02373 5933 5936 5773 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02372 5932 5933 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02371 8185 5932 5772 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02370 5930 5931 5932 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02369 5938 5930 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02368 8185 5930 5938 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02367 7725 7750 7506 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02366 7506 7747 7725 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02365 8185 7793 7506 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02364 4628 4744 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02363 4728 4735 4628 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02362 8185 5453 4047 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02361 4047 8159 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02360 8185 4734 4047 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02359 4030 5670 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02358 4556 4543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02357 6304 5906 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02356 7750 7752 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02355 7766 7247 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02354 8046 7513 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02353 4214 5147 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02352 4213 5148 4214 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02351 8185 7802 4213 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02350 4212 4213 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02349 810 912 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02348 809 914 911 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02347 808 913 907 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02346 8185 1317 808 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02345 8185 1772 913 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02344 914 913 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02343 8185 1074 912 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02342 911 913 810 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02341 909 911 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02340 8185 909 809 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02339 907 914 909 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02338 1317 907 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02337 8185 907 1317 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02336 8185 4995 4250 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02335 7871 4250 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02334 8185 4250 7871 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02333 8185 4250 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02332 8144 4250 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02331 8185 4995 4996 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02330 6383 4996 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02329 8185 4996 6383 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02328 8185 4996 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02327 8144 4996 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02326 8185 4552 4553 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02325 4995 4553 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02324 8185 4553 4995 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02323 8185 4553 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02322 8144 4553 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02321 8185 5616 5617 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02320 5617 6867 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02319 5910 5617 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02318 7527 7791 7526 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02317 7526 7788 7527 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02316 8185 8021 7526 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02315 7525 7527 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02314 4647 7787 2790 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02313 2790 5907 4647 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02312 8185 6792 2790 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02311 1156 2492 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02310 1570 1799 1156 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02309 4009 6273 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02308 4413 6267 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02307 3716 6484 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02306 3602 5180 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02305 4834 5906 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02304 4932 6285 4834 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02303 4833 6286 4932 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02302 8185 5603 4833 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02301 4832 6076 4932 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02300 8185 6284 4832 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02299 4186 1738 1214 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02298 1214 1739 4186 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02297 8185 3148 1214 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02296 3036 3100 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02295 3286 3095 3036 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02294 1203 1296 1202 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02293 1202 2168 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02292 1297 1295 1203 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02291 5233 5236 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02290 5231 5235 5234 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02289 5228 5237 5229 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02288 8185 5227 5228 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02287 8185 5864 5237 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02286 5235 5237 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02285 8185 5232 5236 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02284 5234 5237 5233 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02283 5230 5234 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02282 8185 5230 5231 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02281 5229 5235 5230 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02280 5227 5229 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02279 8185 5229 5227 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02278 6255 6917 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02277 6417 7140 6255 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02276 7683 7871 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02275 8169 8159 7683 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02274 6401 6629 6240 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02273 6240 6400 6401 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02272 8185 6399 6240 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02271 1679 2469 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02270 7550 4572 1679 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02269 1674 5830 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02268 1742 1741 1674 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02267 8185 2177 2065 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02266 2065 4003 2176 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02265 2638 2176 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02264 2060 2166 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02263 2365 3229 2060 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02262 6512 6515 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02261 6511 6514 6510 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02260 6507 6516 6508 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02259 8185 6506 6507 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02258 8185 8063 6516 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02257 6514 6516 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02256 8185 6513 6515 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02255 6510 6516 6512 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02254 6509 6510 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02253 8185 6509 6511 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02252 6508 6514 6509 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02251 6506 6508 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02250 8185 6508 6506 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02249 7066 7352 7067 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02248 7067 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02247 7542 8097 7066 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02246 8185 5574 5575 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02245 5575 5576 5577 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02244 5897 5577 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02243 2926 7314 1265 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02242 8185 1807 1379 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02241 1265 1379 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02240 421 1115 537 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02239 537 1114 422 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02238 422 535 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02237 420 725 537 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02236 8185 1110 420 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02235 8185 739 421 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02234 1965 537 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02233 5793 6300 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02232 5833 5905 5793 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02231 2838 3759 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02230 3114 4166 2838 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02229 8185 5629 5630 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02228 5630 5628 5631 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02227 7747 5631 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02226 5318 5654 5319 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02225 5319 5648 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02224 5317 6796 5318 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02223 5637 6375 5317 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02222 6739 7880 6740 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02221 6740 6909 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02220 6738 6921 6739 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02219 7106 7130 6738 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02218 6641 7398 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02217 6647 7891 6641 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02216 5917 6090 5764 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02215 5764 6089 5917 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02214 8185 6567 5764 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02213 4188 4191 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02212 6466 4186 4188 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02211 1710 2132 1632 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02210 1632 3737 1710 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02209 8185 2599 1632 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02208 2802 3566 2804 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02207 2804 3293 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02206 2801 3586 2802 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02205 2803 3581 2801 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02204 8185 3556 2859 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02203 2858 3135 2852 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02202 2856 3129 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_02201 2852 2854 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02200 8185 3556 2854 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_02199 2860 2858 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_02198 2859 2853 2855 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02197 2855 3129 2858 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02196 2858 2856 2857 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02195 2857 3145 2859 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02194 8185 3556 2538 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02193 2656 2648 2536 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02192 2650 3129 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_02191 2536 2651 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02190 8185 3556 2651 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_02189 2873 2656 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_02188 2538 2652 2537 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02187 2537 3129 2656 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02186 2656 2650 2539 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02185 2539 3143 2538 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_02184 6216 6307 6217 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02183 6217 6309 6310 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02182 8185 6308 6216 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02181 6536 6310 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_02180 8185 7343 4718 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02179 4718 4720 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02178 5437 4719 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02177 4718 4717 4719 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02176 4719 6363 4718 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02175 7092 7867 7091 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02174 8185 7091 7884 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02173 8185 7867 7094 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02172 7093 7549 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02171 7091 7094 7093 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02170 8185 7272 7092 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_02169 7884 7091 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02168 5308 5618 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_02167 5616 5620 5308 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_02166 5307 5428 5616 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_02165 8185 5429 5307 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_02164 5307 5432 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_02163 1538 5624 1537 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02162 1537 4293 1538 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02161 8185 1992 1537 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02160 8185 8179 5787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02159 5787 5971 5970 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02158 6178 5970 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02157 8185 4251 4252 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02156 4252 7871 4253 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02155 4756 4253 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02154 5255 7633 5254 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02153 5254 6909 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02152 5253 6172 5255 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02151 5503 7130 5253 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02150 7757 7758 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02149 8185 7787 7757 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02148 7757 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02147 8185 8045 7757 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02146 8004 7757 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02145 2563 5434 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02144 8185 2698 2563 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02143 2563 4548 2700 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02142 2700 2702 2563 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02141 5744 7314 7073 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02140 8185 7314 5881 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02139 5743 5888 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02138 7073 5881 5743 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02137 8185 5880 5744 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02136 3344 4517 3347 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02135 3347 4228 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02134 3345 7343 3344 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02133 3583 4518 3345 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02132 3232 5648 3233 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02131 3233 6543 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02130 3231 6544 3232 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02129 3320 3322 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02128 3322 6267 3231 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02127 4416 4914 4335 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02126 4335 4502 4416 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02125 8185 4503 4335 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02124 8185 6172 6173 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02123 6173 6909 6175 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02122 6407 6175 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02121 8185 5089 4819 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02120 4819 5566 4899 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02119 4898 4899 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02118 8185 342 35 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02117 35 343 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02116 1115 156 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02115 35 159 156 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02114 156 163 35 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02113 4224 4538 4222 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02112 8185 4720 4223 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02111 4222 4223 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02110 8185 7352 5364 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02109 5364 5718 5506 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02108 5505 5506 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02107 8185 3244 3028 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02106 3028 3156 3157 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02105 3165 3157 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02104 8185 1541 1121 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02103 1121 1119 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02102 1785 1122 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02101 1121 1535 1122 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02100 1122 1120 1121 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_02099 6482 6484 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02098 6483 6480 6482 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02097 8185 6481 6483 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02096 6478 6483 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02095 6193 6267 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02094 6265 6480 6193 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02093 8185 6266 6265 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02092 6661 7884 6662 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02091 6662 7892 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02090 6659 6893 6661 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02089 6658 6660 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02088 6660 7891 6659 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02087 5084 5087 5384 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02086 8185 5938 5084 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02085 5086 5453 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02084 5384 5085 5086 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02083 8185 5453 5087 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02082 5085 5938 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02081 4045 8064 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02080 8185 5863 4045 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02079 2580 6797 2581 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02078 2581 6802 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02077 2579 4302 2580 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02076 2951 2721 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_02075 2721 3857 2579 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02074 2998 3763 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02073 3127 4424 2998 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02072 8185 4510 3127 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02071 414 524 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02070 413 525 523 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02069 412 526 519 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02068 8185 517 412 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02067 8185 1772 526 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02066 525 526 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02065 8185 528 524 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02064 523 526 414 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02063 521 523 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02062 8185 521 413 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02061 519 525 521 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02060 517 519 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02059 8185 519 517 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02058 6228 6371 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02057 6229 6372 6369 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02056 6227 6373 6366 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02055 8185 6602 6227 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02054 8185 7821 6373 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02053 6372 6373 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02052 8185 6600 6371 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02051 6369 6373 6228 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02050 6367 6369 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02049 8185 6367 6229 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02048 6366 6372 6367 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02047 6602 6366 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02046 8185 6366 6602 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02045 5747 5891 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02044 5748 5892 5890 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02043 5746 5893 5887 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02042 8185 5888 5746 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02041 8185 8063 5893 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02040 5892 5893 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02039 8185 7528 5891 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02038 5890 5893 5747 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02037 5889 5890 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02036 8185 5889 5748 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02035 5887 5892 5889 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02034 5888 5887 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02033 8185 5887 5888 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02032 8185 7789 8028 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02031 8028 7782 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02030 8185 7783 8028 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02029 4074 4070 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02028 8185 4315 4074 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02027 4074 4071 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02026 8185 4472 4074 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02025 9 79 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02024 8 80 76 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02023 7 81 73 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02022 8185 498 7 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02021 8185 1951 81 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02020 80 81 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_02019 8185 261 79 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_02018 76 81 9 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02017 75 76 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02016 8185 75 8 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02015 73 80 75 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02014 498 73 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02013 8185 73 498 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_02012 8185 7257 7460 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02011 7460 6820 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02010 8185 6816 7460 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02009 1473 1739 1209 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02008 1209 1738 1473 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02007 8185 8045 1209 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02006 3659 3667 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02005 8185 3656 3659 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02004 3659 3851 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02003 8185 4078 3659 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_02002 3802 3801 3803 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02001 3803 4033 3802 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_02000 8185 3804 3803 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01999 4856 5010 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01998 4855 5011 5009 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01997 4854 5012 5005 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01996 8185 5003 4854 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01995 8185 5864 5012 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01994 5011 5012 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01993 8185 5226 5010 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01992 5009 5012 4856 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01991 5006 5009 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01990 8185 5006 4855 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01989 5005 5011 5006 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01988 5003 5005 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01987 8185 5005 5003 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01986 1630 1707 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01985 1631 1706 1704 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01984 1629 1708 1701 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01983 8185 5453 1629 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01982 8185 3708 1708 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01981 1706 1708 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01980 8185 2319 1707 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01979 1704 1708 1630 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01978 1702 1704 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01977 8185 1702 1631 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01976 1701 1706 1702 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01975 5453 1701 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01974 8185 1701 5453 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01973 7222 7309 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01972 7310 7314 7222 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01971 7661 7772 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01970 8038 7773 7661 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01969 5736 5875 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01968 6188 6672 5736 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01967 7225 7321 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01966 7458 7322 7225 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01965 3336 3581 3337 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01964 3337 3356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01963 3553 3582 3336 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01962 1457 2796 1456 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01961 1456 3744 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01960 1455 3542 1457 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01959 2159 1739 1646 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01958 1646 1738 2159 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01957 8185 1962 1646 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01956 5611 5614 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01955 5610 5613 5612 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01954 5607 5615 5608 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01953 8185 5606 5607 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01952 8185 8063 5615 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01951 5613 5615 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01950 8185 5846 5614 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01949 5612 5615 5611 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01948 5609 5612 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01947 8185 5609 5610 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01946 5608 5613 5609 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01945 5606 5608 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01944 8185 5608 5606 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01943 4227 4310 4226 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01942 4226 4224 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01941 4225 6609 4227 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01940 5161 6796 4225 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01939 6165 6652 6167 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01938 6167 7121 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01937 6166 6636 6165 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01936 3015 4302 3014 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01935 3014 6609 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01934 5908 5654 3015 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01933 3852 3850 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01932 3851 4287 3852 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01931 2221 2896 2095 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01930 2094 6796 2221 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01929 2095 4067 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01928 2220 2221 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01927 8185 2894 2094 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01926 2094 2688 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01925 2348 3730 2347 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01924 2347 3735 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01923 2346 3348 2348 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01922 2668 2661 2543 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01921 2543 2659 2668 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01920 8185 2883 2543 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01919 4815 4892 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01918 4816 4893 4890 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01917 4814 4894 4887 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01916 8185 6349 4814 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01915 8185 8063 4894 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01914 4893 4894 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01913 8185 5090 4892 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01912 4890 4894 4815 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01911 4888 4890 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01910 8185 4888 4816 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01909 4887 4893 4888 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01908 6349 4887 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01907 8185 4887 6349 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01906 8185 7523 7521 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01905 7521 7520 7522 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01904 7748 7522 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01903 4850 5000 4851 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01902 4851 4997 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01901 4998 4999 4850 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01900 5714 5870 5713 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01899 5713 6404 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01898 5712 5728 5714 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01897 6243 6663 6244 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01896 6244 6642 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01895 6404 7887 6243 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01894 3627 6598 3491 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01893 3491 3625 3627 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01892 8185 3628 3491 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01891 3624 3627 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01890 3786 3794 3785 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01889 3785 3788 3784 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01888 8185 4203 3786 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01887 3783 3784 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01886 8185 3566 2510 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01885 2510 3293 2604 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01884 2602 2604 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01883 3736 4172 3734 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01882 3734 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01881 3735 7585 3736 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01880 655 6867 656 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01879 8185 656 654 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01878 8185 6867 658 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01877 657 3276 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01876 656 658 657 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01875 8185 6520 655 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01874 654 656 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01873 4643 6867 4642 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01872 8185 4642 4641 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01871 8185 6867 4645 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01870 4646 4644 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01869 4642 4645 4646 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01868 8185 6292 4643 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01867 4641 4642 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01866 3880 6867 3960 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01865 8185 3960 3955 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01864 8185 6867 3961 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01863 3881 3958 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01862 3960 3961 3881 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01861 8185 3956 3880 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01860 3955 3960 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01859 3381 3378 3380 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01858 3380 3618 3383 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01857 8185 3379 3381 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01856 5426 3383 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01855 5352 7633 5353 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01854 5353 5971 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01853 5498 5868 5352 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01852 3170 1800 1663 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01851 1663 1798 3170 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01850 8185 3150 1663 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01849 348 1150 350 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01848 350 359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01847 349 4558 348 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01846 3882 6867 3966 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01845 8185 3966 3962 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01844 8185 6867 3967 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01843 3883 3964 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01842 3966 3967 3883 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01841 8185 6792 3882 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01840 3962 3966 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01839 5762 7026 5761 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01838 5761 6543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01837 5760 7353 5762 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01836 6554 6080 5760 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01835 7564 7957 7591 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01834 8185 7957 7563 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01833 7565 7835 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01832 7591 7563 7565 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01831 8185 7970 7564 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01830 4813 5880 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01829 5373 7500 4813 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01828 7771 8009 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01827 8185 7787 7771 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01826 7771 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01825 8185 8045 7771 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01824 7773 7771 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01823 5089 7787 5088 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01822 5088 5907 5089 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01821 8185 6349 5088 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01820 8185 4734 3837 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01819 8185 8159 3837 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01818 3837 5453 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01817 3839 3837 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01816 6195 6485 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01815 6270 7500 6195 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01814 8185 4953 4342 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01813 4342 4932 4513 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01812 4427 4513 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01811 7234 7408 7235 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01810 7235 7881 7394 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01809 8185 7883 7234 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01808 7872 7394 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01807 8185 3714 3712 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01806 3712 4130 3713 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01805 3711 3713 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01804 3724 4413 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01803 8185 7787 3724 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01802 3724 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01801 8185 8045 3724 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01800 3723 3724 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01799 7063 7957 7612 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01798 8185 7957 7065 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01797 7064 7558 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01796 7612 7065 7064 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01795 8185 7803 7063 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01794 8185 5148 3779 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01793 3779 5147 3778 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01792 3776 3778 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01791 8185 166 44 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01790 44 365 162 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01789 161 162 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01788 1954 4189 1955 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01787 1955 2170 1954 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01786 8185 2375 1955 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01785 6644 7892 6643 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01784 6643 7398 6645 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01783 8185 7869 6644 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01782 6642 6645 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01781 4817 4902 4818 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01780 4818 4896 4897 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01779 8185 5606 4817 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01778 4895 4897 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01777 1686 7051 1687 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01776 1687 2719 1828 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01775 8185 3857 1686 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01774 1827 1828 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01773 6246 6893 6245 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01772 6245 7881 6405 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01771 8185 7891 6246 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01770 6636 6405 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01769 17 101 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01768 16 103 100 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01767 15 104 96 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01766 8185 273 15 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01765 8185 1951 104 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01764 103 104 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01763 8185 272 101 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01762 100 104 17 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01761 99 100 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01760 8185 99 16 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01759 96 103 99 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01758 273 96 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01757 8185 96 273 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01756 7311 7247 6677 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01755 8185 7957 6762 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01754 6677 6762 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01753 3813 4302 3814 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01752 3814 4068 3815 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01751 8185 4574 3813 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01750 3812 3815 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01749 837 6802 838 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01748 838 4575 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01747 836 4068 837 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01746 1167 958 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01745 958 6796 836 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01744 5417 6506 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01743 4406 6489 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01742 4705 6775 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01741 2361 1956 1494 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01740 1494 1957 2361 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01739 8185 1962 1494 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01738 2835 3111 2834 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01737 2834 3112 2835 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01736 8185 3108 2834 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01735 2833 2835 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01734 5335 5475 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01733 5334 5477 5474 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01732 5333 5476 5470 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01731 8185 5664 5333 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01730 8185 5864 5476 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01729 5477 5476 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01728 8185 5478 5475 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01727 5474 5476 5335 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01726 5471 5474 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01725 8185 5471 5334 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01724 5470 5477 5471 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01723 5664 5470 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01722 8185 5470 5664 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01721 5288 7352 5289 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01720 5289 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01719 5896 5394 5288 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01718 5111 5118 5112 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01717 5112 5113 5111 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01716 8185 5110 5112 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01715 5109 5111 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01714 3249 3623 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01713 3252 4048 3249 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01712 4999 5202 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01711 6594 6602 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01710 4260 5227 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01709 4032 4760 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01708 5429 5603 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01707 5413 5898 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01706 1503 1508 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01705 1505 1507 1504 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01704 1500 1509 1501 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01703 8185 1499 1500 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01702 8185 1772 1509 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01701 1507 1509 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01700 8185 1506 1508 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01699 1504 1509 1503 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01698 1502 1504 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01697 8185 1502 1505 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01696 1501 1507 1502 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01695 1499 1501 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01694 8185 1501 1499 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01693 4265 4268 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01692 4264 4267 4266 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01691 4261 4269 4262 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01690 8185 4770 4261 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01689 8185 5864 4269 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01688 4267 4269 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01687 8185 4769 4268 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01686 4266 4269 4265 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01685 4263 4266 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01684 8185 4263 4264 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01683 4262 4267 4263 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01682 4770 4262 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01681 8185 4262 4770 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01680 8033 8036 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01679 8032 8035 8034 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01678 8029 8037 8030 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01677 8185 8040 8029 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01676 8185 8063 8037 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01675 8035 8037 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01674 8185 8039 8036 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01673 8034 8037 8033 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01672 8031 8034 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01671 8185 8031 8032 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01670 8030 8035 8031 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01669 8040 8030 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01668 8185 8030 8040 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01667 5301 7352 5300 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01666 5300 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01665 6298 5419 5301 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01664 1680 7356 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01663 1798 5942 1680 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01662 6524 6292 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01661 2035 1389 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01660 8185 1390 2035 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01659 2035 1615 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01658 8185 1616 2035 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01657 2063 4427 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01656 2502 2172 2063 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01655 7309 7318 7166 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01654 7166 7503 7309 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01653 8185 7316 7166 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01652 827 3608 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01651 956 957 827 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01650 952 946 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01649 8185 947 952 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01648 952 1139 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01647 8185 948 952 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01646 1119 952 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01645 5240 5502 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01644 5241 5724 5240 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01643 5797 5944 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01642 6128 6137 5797 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01641 5663 5937 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01640 5944 6127 5663 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01639 7689 7881 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01638 7882 7891 7689 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01637 7646 7643 7644 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01636 7644 8186 7646 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01635 8185 7869 7644 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01634 2719 5940 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01633 8185 2262 2719 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01632 2719 2964 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01631 8185 2968 2719 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01630 8185 5197 3458 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01629 3458 3780 3580 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01628 3579 3580 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01627 5584 5583 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01626 5581 5585 5582 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01625 5578 5586 5579 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01624 8185 5898 5578 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01623 8185 8063 5586 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01622 5585 5586 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01621 8185 5589 5583 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01620 5582 5586 5584 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01619 5580 5582 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01618 8185 5580 5581 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01617 5579 5585 5580 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01616 5898 5579 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01615 8185 5579 5898 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01614 6082 7352 6081 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01613 6081 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01612 6309 6080 6082 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01611 8185 5665 5332 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01610 5332 5682 5468 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01609 5467 5468 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01608 7196 8140 7371 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01607 8185 7371 7271 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01606 8185 8140 7275 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01605 7197 7549 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01604 7371 7275 7197 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01603 8185 7272 7196 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01602 7271 7371 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01601 7198 8140 7375 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01600 8185 7375 7575 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01599 8185 8140 7278 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01598 7199 7528 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01597 7375 7278 7199 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01596 8185 7572 7198 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01595 7575 7375 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01594 7577 8140 7579 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01593 8185 7579 7851 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01592 8185 8140 7580 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01591 7578 7585 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01590 7579 7580 7578 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01589 8185 7845 7577 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01588 7851 7579 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01587 7206 8140 7386 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01586 8185 7386 7384 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01585 8185 8140 7289 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01584 7207 7349 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01583 7386 7289 7207 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01582 8185 7379 7206 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01581 7384 7386 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01580 7605 8140 7606 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01579 8185 7606 7603 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01578 8185 8140 7608 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01577 7607 7777 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01576 7606 7608 7607 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01575 8185 7604 7605 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01574 7603 7606 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01573 6714 7867 6852 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01572 8185 6852 6907 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01571 8185 7867 6853 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01570 6715 6850 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01569 6852 6853 6715 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01568 8185 7076 6714 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01567 6907 6852 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01566 3437 4574 3436 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01565 3436 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01564 3435 7353 3437 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01563 3542 6484 3435 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01562 8138 8140 8142 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01561 8185 8142 8153 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01560 8185 8140 8143 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01559 8141 8139 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01558 8142 8143 8141 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01557 8185 8147 8138 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01556 8153 8142 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01555 7598 8140 7861 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01554 8185 7861 8130 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01553 8185 8140 7862 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01552 7602 7863 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01551 7861 7862 7602 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01550 8185 8125 7598 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01549 8130 7861 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01548 5490 6629 5343 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01547 5343 5866 5490 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01546 8185 5489 5343 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01545 4309 4575 4308 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01544 4308 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01543 4307 4306 4309 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01542 4317 5483 4307 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01541 7322 7797 7172 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01540 7172 7798 7322 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01539 8185 7528 7172 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01538 1472 1943 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01537 1936 2154 1472 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01536 8185 2616 1936 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01535 3452 4167 3451 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01534 3451 6543 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01533 3450 6544 3452 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01532 3566 6267 3450 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01531 4709 5434 4708 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01530 4708 5574 4710 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01529 8185 6363 4709 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01528 4707 4710 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01527 2077 2203 2078 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01526 2078 7343 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01525 2076 5148 2077 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01524 4172 2204 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01523 2204 4548 2076 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01522 5672 6383 5673 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01521 8185 5673 5671 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01520 8185 6383 5675 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01519 5674 5858 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01518 5673 5675 5674 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01517 8185 5670 5672 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01516 5671 5673 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01515 7597 7867 7600 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01514 8185 7600 7643 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01513 8185 7867 7601 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01512 7599 7863 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01511 7600 7601 7599 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01510 8185 8125 7597 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01509 7643 7600 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01508 1677 1788 1678 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01507 1678 2214 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01506 1676 1985 1677 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01505 4173 1789 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01504 1789 2207 1676 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01503 6502 6784 6204 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01502 6204 6785 6502 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01501 8185 7500 6204 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01500 7400 7304 7152 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01499 7152 7151 7400 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01498 8185 7149 7152 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01497 6160 6156 6159 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01496 6159 6157 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01495 6155 6158 6160 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01494 6154 6166 6155 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01493 4699 4696 4698 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01492 8185 7059 4699 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01491 4700 5120 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01490 4698 4697 4700 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01489 8185 5120 4696 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01488 4697 7059 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01487 6765 6972 6679 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01486 6678 7550 6765 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01485 6679 6985 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01484 6763 6765 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01483 8185 7548 6678 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01482 6678 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01481 4490 4406 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01480 8185 7787 4490 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01479 4490 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01478 8185 8045 4490 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01477 4405 4490 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01476 1315 1956 1217 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01475 1217 1957 1315 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01474 8185 8045 1217 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01473 1673 1818 1672 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01472 1672 1817 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01471 1671 1816 1673 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01470 2466 1819 1671 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01469 1313 1957 1215 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01468 1215 1956 1313 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01467 8185 3148 1215 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01466 796 860 3276 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01465 8185 2595 796 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01464 797 865 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01463 3276 858 797 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01462 8185 865 860 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01461 858 2595 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01460 7518 8046 7519 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01459 7519 7747 7518 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01458 8185 7517 7519 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01457 7549 6850 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01456 8185 4790 3947 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01455 3947 5032 4066 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01454 4071 4066 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01453 8185 1335 1224 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01452 1224 5641 1329 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01451 1327 1329 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01450 4183 7056 4182 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01449 4182 5406 4183 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01448 8185 6812 4182 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01447 6780 6781 6684 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01446 6684 6778 6780 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01445 8185 6779 6684 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01444 5809 8187 5808 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01443 5808 7881 5969 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01442 8185 7883 5809 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01441 5971 5969 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01440 8185 5483 767 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01439 767 4310 769 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01438 1140 769 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01437 2103 2235 2102 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01436 2102 2234 2237 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01435 8185 2236 2103 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01434 2246 2237 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01433 6325 6375 5769 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01432 5769 5922 6325 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01431 8185 5923 5769 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01430 4805 4802 4804 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01429 4804 4803 4806 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01428 8185 5044 4805 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01427 4801 4806 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01426 1756 1964 1651 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01425 1651 1965 1756 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01424 8185 1962 1651 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01423 2174 1756 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01422 3128 2178 1963 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01421 1963 2179 3128 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01420 8185 1962 1963 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01419 28 138 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01418 29 139 137 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01417 27 140 133 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01416 8185 530 27 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01415 8185 1772 140 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01414 139 140 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01413 8185 141 138 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01412 137 140 28 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01411 134 137 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01410 8185 134 29 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01409 133 139 134 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01408 530 133 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01407 8185 133 530 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01406 361 558 362 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01405 362 559 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01404 360 1362 361 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01403 359 358 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01402 358 6363 360 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01401 706 1115 708 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01400 708 1114 707 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01399 707 709 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01398 705 703 708 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01397 8185 1110 705 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01396 8185 900 706 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01395 1957 708 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01394 1118 1113 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01393 1348 1114 1118 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01392 1117 1115 1348 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01391 8185 1116 1117 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01390 1112 1111 1348 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01389 8185 1110 1112 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01388 1930 2138 1931 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01387 1931 2595 1930 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01386 8185 1929 1931 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01385 1928 1930 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01384 60 197 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01383 59 198 196 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01382 58 199 192 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01381 8185 190 58 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01380 8185 3834 199 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01379 198 199 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01378 8185 1699 197 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01377 196 199 60 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01376 193 196 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01375 8185 193 59 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01374 192 198 193 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01373 190 192 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01372 8185 192 190 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01371 6980 6981 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01370 6978 6982 6979 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01369 6975 6983 6976 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01368 8185 6974 6975 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01367 8185 8063 6983 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01366 6982 6983 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01365 8185 7585 6981 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01364 6979 6983 6980 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01363 6977 6979 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01362 8185 6977 6978 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01361 6976 6982 6977 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01360 6974 6976 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01359 8185 6976 6974 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01358 8185 8053 8067 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01357 8067 8054 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01356 8185 8052 8067 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01355 7359 7056 7057 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01354 7057 7058 7359 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01353 8185 7342 7057 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01352 1270 4295 1271 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01351 1271 4310 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01350 1269 4167 1270 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01349 1384 1385 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01348 1385 5624 1269 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01347 3611 4032 3472 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01346 3472 3610 3611 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01345 8185 3613 3472 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01344 750 753 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01343 643 752 748 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01342 642 754 747 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01341 8185 1116 642 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01340 8185 3834 754 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01339 752 754 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01338 8185 751 753 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01337 748 754 750 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01336 749 748 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01335 8185 749 643 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01334 747 752 749 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01333 1116 747 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01332 8185 747 1116 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01331 6623 6626 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01330 6621 6625 6624 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01329 6619 6628 6620 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01328 8185 6618 6619 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01327 8185 8166 6628 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01326 6625 6628 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01325 8185 6630 6626 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01324 6624 6628 6623 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01323 6622 6624 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01322 8185 6622 6621 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01321 6620 6625 6622 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01320 6618 6620 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01319 8185 6620 6618 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01318 4246 4247 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01317 4243 4248 4245 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01316 4240 4249 4241 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01315 8185 4955 4240 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01314 8185 5864 4249 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01313 4248 4249 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01312 8185 4244 4247 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01311 4245 4249 4246 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01310 4242 4245 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01309 8185 4242 4243 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01308 4241 4248 4242 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01307 4955 4241 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01306 8185 4241 4955 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01305 242 3956 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01304 8185 3956 241 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01303 8185 2127 239 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01302 240 238 242 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01301 239 241 240 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01300 1446 240 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01299 8185 240 1446 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01298 238 2127 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01297 6253 6921 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01296 6412 7148 6253 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01295 6252 7151 6412 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01294 8185 6655 6252 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01293 6252 6658 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01292 8026 8028 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01291 8066 8025 8026 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01290 7556 7791 7555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01289 7555 7788 7556 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01288 8185 8071 7555 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01287 8053 7556 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01286 2316 2789 2317 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01285 2317 5633 2316 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01284 8185 5372 2317 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01283 2315 2316 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01282 4578 4583 4374 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01281 4374 5245 4578 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01280 8185 4577 4374 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01279 4468 4578 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01278 3462 3794 3463 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01277 3463 3788 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01276 3587 4203 3462 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01275 3339 3579 3338 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01274 3338 3356 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01273 3737 3582 3339 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01272 2045 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01271 2133 2135 2045 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01270 2044 2599 2133 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01269 8185 2132 2044 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01268 2044 3737 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_01267 794 855 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01266 795 856 853 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01265 793 857 850 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01264 8185 2127 793 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01263 8185 3708 857 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01262 856 857 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01261 8185 2126 855 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01260 853 857 794 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01259 851 853 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01258 8185 851 795 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01257 850 856 851 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01256 2127 850 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01255 8185 850 2127 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01254 7145 7884 7146 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01253 7146 7403 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01252 7147 8184 7145 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01251 7461 7460 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01250 8089 7801 7461 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01249 3954 4474 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01248 4078 4477 3954 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01247 2029 2251 2028 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01246 2028 2448 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01245 2242 2027 2029 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01244 4843 4965 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01243 4842 4967 4961 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01242 4841 4966 4958 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01241 8185 6341 4841 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01240 8185 7821 4966 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01239 4967 4966 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01238 8185 4963 4965 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01237 4961 4966 4843 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01236 4960 4961 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01235 8185 4960 4842 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01234 4958 4967 4960 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01233 6341 4958 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01232 8185 4958 6341 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01231 4824 4910 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01230 4823 4911 4909 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01229 4822 4912 4905 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01228 8185 6801 4822 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01227 8185 8063 4912 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01226 4911 4912 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_01225 8185 4913 4910 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01224 4909 4912 4824 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01223 4906 4909 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01222 8185 4906 4823 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01221 4905 4911 4906 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01220 6801 4905 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01219 8185 4905 6801 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01218 6266 6793 5554 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01217 5554 6294 6266 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01216 8185 5553 5554 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01215 8185 5160 5163 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01214 5163 5161 5165 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01213 5162 5165 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01212 8094 1790 1660 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01211 1660 1785 8094 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01210 8185 7314 1660 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01209 6470 7738 6471 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01208 6471 7730 6470 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01207 8185 8064 6471 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01206 6469 6470 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01205 8185 6341 3467 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01204 3467 3611 3604 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01203 3603 3604 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01202 1466 1476 1207 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01201 1207 1477 1466 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01200 8185 1962 1207 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01199 8185 7012 5125 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01198 5125 5164 5126 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01197 5124 5126 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01196 4675 6867 4917 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01195 8185 4917 4913 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01194 8185 6867 4918 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01193 4678 4914 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01192 4917 4918 4678 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01191 8185 6801 4675 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01190 4913 4917 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01189 5091 6867 5094 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01188 8185 5094 5090 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01187 8185 6867 5095 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01186 5093 5092 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01185 5094 5095 5093 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01184 8185 6349 5091 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01183 5090 5094 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01182 6048 6500 6049 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01181 6049 6051 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01180 6047 6786 6048 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01179 6262 6503 6047 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01178 5784 6921 5785 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01177 5785 6909 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01176 5870 5968 5784 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01175 759 5483 758 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01174 758 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01173 760 1353 759 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01172 8185 2202 1775 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01171 1775 2199 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01170 1776 1775 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01169 4336 6867 4509 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01168 8185 4509 4681 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01167 8185 6867 4423 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01166 4337 4502 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01165 4509 4423 4337 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01164 8185 6549 4336 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_01163 4681 4509 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01162 7545 7541 7544 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01161 7544 7542 7546 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01160 8185 7543 7545 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01159 7794 7546 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01158 4117 6472 4119 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01157 4119 6478 4118 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01156 8185 6473 4117 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01155 5078 4118 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01154 6201 6786 6202 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01153 6202 6500 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01152 6200 6784 6201 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01151 6778 6281 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01150 6281 6785 6200 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01149 6335 6618 6017 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01148 8185 6549 6018 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01147 6017 6018 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01146 7215 7300 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01145 7395 7875 7215 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01144 8185 7871 7395 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01143 7297 7395 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01142 8185 7405 6669 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01141 6669 6670 6671 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01140 6668 6671 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01139 5727 5875 5729 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01138 5729 6176 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01137 5728 6921 5727 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01136 8185 1807 1160 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01135 1160 8064 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01134 2698 1160 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01133 8185 8159 2923 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01132 2923 5453 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01131 2922 2923 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01130 8185 5940 2261 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01129 2122 2261 2260 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01128 8185 2262 2122 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01127 2490 2260 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01126 8185 2260 2490 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01125 6529 6804 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01124 6532 7500 6529 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01123 1987 7548 1988 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01122 1988 7559 1987 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01121 8185 1986 1988 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01120 2205 1987 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01119 1453 2135 1454 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01118 1452 2599 1453 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01117 1454 3744 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01116 1451 1453 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01115 8185 2132 1452 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01114 1452 3737 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_01113 3728 4167 3729 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01112 3729 6797 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01111 3726 6796 3728 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01110 3725 3727 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01109 3727 6273 3726 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01108 6540 7797 6539 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01107 6539 7798 6540 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01106 8185 8122 6539 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01105 8185 5967 5783 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01104 5783 6409 5966 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01103 5869 5966 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01102 8049 8046 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01101 8185 8047 8049 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01100 8049 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01099 8185 8045 8049 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01098 8068 8049 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01097 4376 6672 4377 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01096 4377 6421 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01095 4375 4790 4376 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01094 4470 5740 4375 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01093 6973 6987 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01092 6972 7957 6973 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01091 1886 6359 1888 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01090 1888 1887 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01089 1885 2924 1886 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01088 2207 1994 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01087 1994 1891 1885 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01086 7459 6793 6692 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01085 6692 7058 7459 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01084 8185 6794 6692 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01083 8185 5913 5759 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01082 5759 5912 5914 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01081 5837 5914 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01080 7667 7803 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01079 7804 7957 7667 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01078 5973 7893 5788 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01077 5788 7408 5973 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01076 8185 8184 5788 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01075 5876 5973 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01074 8185 4801 4800 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01073 4800 5034 4799 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01072 4798 4799 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01071 8185 4318 3878 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01070 3878 3877 3879 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01069 3876 3879 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01068 8185 2227 2081 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01067 2081 7343 2208 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01066 2421 2208 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01065 4341 4511 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01064 4426 4512 4341 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01063 8185 4510 4426 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01062 6744 7884 6745 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01061 6745 7403 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01060 6743 7408 6744 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01059 6917 6911 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01058 6911 8184 6743 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01057 8185 1304 1210 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01056 1210 5641 1305 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01055 1739 1305 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01054 2341 2614 2342 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01053 2342 3725 2341 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01052 8185 3315 2342 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01051 2340 2341 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01050 7488 7486 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01049 7487 7490 7488 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01048 8185 7484 7487 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01047 7485 7487 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01046 3398 4573 3400 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01045 3400 6311 3401 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01044 8185 4293 3398 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01043 3844 3401 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01042 3263 3260 3265 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01041 3265 3659 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01040 3262 3858 3263 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01039 3419 3418 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01038 3418 3261 3262 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01037 3047 4203 3048 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01036 3048 3794 3149 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01035 8185 5908 3047 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01034 3148 3149 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01033 8185 7314 1450 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01032 1449 1450 1448 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01031 8185 6267 1449 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01030 6084 1448 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01029 8185 1448 6084 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_01028 8185 6870 6607 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01027 6607 7095 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01026 8185 6618 6607 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01025 3474 4306 3473 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01024 3473 6609 3617 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01023 8185 5447 3474 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01022 3809 3617 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01021 3055 3182 3056 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01020 3056 3416 3181 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01019 8185 3410 3055 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01018 3187 3181 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_01017 2120 4293 2121 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01016 2121 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01015 2119 5648 2120 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01014 2258 2259 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01013 2259 5654 2119 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01012 5259 5265 5260 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01011 5260 5505 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01010 5257 5730 5259 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01009 5256 5258 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01008 5258 5262 5257 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01007 4877 6185 4878 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01006 4878 5040 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01005 4876 5256 4877 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01004 5034 5035 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_01003 5035 5036 4876 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_01002 689 693 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_01001 635 692 686 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_01000 634 694 684 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00999 8185 685 634 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00998 8185 1951 694 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00997 692 694 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00996 8185 691 693 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00995 686 694 689 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00994 688 686 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00993 8185 688 635 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00992 684 692 688 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00991 685 684 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00990 8185 684 685 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00989 3932 4041 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00988 3933 4042 4039 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00987 3931 4043 4036 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00986 8185 4255 3931 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00985 8185 5864 4043 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00984 4042 4043 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00983 8185 4254 4041 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00982 4039 4043 3932 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00981 4037 4039 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00980 8185 4037 3933 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00979 4036 4042 4037 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00978 4255 4036 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00977 8185 4036 4255 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00976 6793 6520 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00975 4896 5453 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00974 7020 6792 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00973 6821 6541 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00972 7029 6349 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00971 7056 6801 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00970 3184 2252 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00969 8185 2254 3184 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00968 8185 4688 3758 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00967 3758 3997 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00966 3757 3758 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00965 3119 3121 2996 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00964 2996 3575 3119 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00963 8185 3118 2996 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00962 3310 3119 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00961 720 721 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00960 637 722 716 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00959 636 723 715 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00958 8185 1088 636 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00957 8185 1772 723 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00956 722 723 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00955 8185 915 721 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00954 716 723 720 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00953 718 716 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00952 8185 718 637 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00951 715 722 718 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00950 1088 715 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00949 8185 715 1088 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00948 5573 7041 5572 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00947 5572 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00946 5576 5571 5573 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00945 4717 4538 4348 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00944 4348 4530 4717 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00943 8185 5443 4348 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00942 5794 5908 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00941 5842 6363 5794 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00940 7531 7779 7530 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00939 7530 7778 7531 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00938 8185 7528 7530 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00937 7529 7531 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00936 2099 2235 2098 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00935 2098 2234 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00934 2241 2236 2099 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00933 2247 1173 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00932 8185 1167 2247 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00931 2247 1168 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00930 8185 1169 2247 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00929 2914 2912 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00928 3251 2913 2914 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00927 4901 5108 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00926 4902 5938 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00925 7059 6549 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00924 4939 6076 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00923 2484 1898 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00922 8185 2454 2484 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00921 2484 1897 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00920 8185 2249 2484 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00919 2047 2591 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00918 2594 2143 2047 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00917 8081 8082 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00916 8080 8083 8079 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00915 8076 8084 8077 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00914 8185 8086 8076 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00913 8185 8166 8084 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00912 8083 8084 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00911 8185 8085 8082 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00910 8079 8084 8081 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00909 8078 8079 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00908 8185 8078 8080 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00907 8077 8083 8078 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00906 8086 8077 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00905 8185 8077 8086 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00904 1236 1352 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00903 1539 1353 1236 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00902 1235 2210 1539 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00901 8185 5624 1235 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00900 1235 4293 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00899 5796 6132 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00898 5935 5939 5796 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00897 3919 7354 3918 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00896 3918 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00895 4525 6293 3919 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00894 3817 6311 3816 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00893 3816 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00892 4540 6293 3817 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00891 1253 4068 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00890 1571 4574 1253 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00889 2685 2687 2554 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00888 2553 3370 2685 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00887 2554 2688 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00886 7778 2685 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00885 8185 4067 2553 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00884 2553 4293 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00883 8185 2361 1947 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00882 1947 4685 1949 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00881 2352 1949 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00880 5596 5598 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00879 5595 5597 5594 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00878 5591 5599 5592 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00877 8185 5603 5591 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00876 8185 8063 5599 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00875 5597 5599 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00874 8185 5835 5598 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00873 5594 5599 5596 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00872 5593 5594 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00871 8185 5593 5595 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00870 5592 5597 5593 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00869 5603 5592 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00868 8185 5592 5603 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00867 8185 7343 6074 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00866 6074 6554 6075 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00865 6308 6075 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00864 8185 7343 5560 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00863 5560 5562 5561 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00862 5886 5561 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00861 8120 8140 8121 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00860 8185 8121 8118 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00859 8185 8140 8124 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00858 8123 8122 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00857 8121 8124 8123 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00856 8185 8119 8120 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00855 8118 8121 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00854 5795 5937 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00853 5939 5938 5795 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00852 441 6609 440 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00851 440 1565 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00850 2203 4302 441 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00849 1256 6802 1255 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00848 1255 1565 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00847 2227 4302 1256 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00846 5905 1744 1647 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00845 1647 1743 5905 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00844 8185 3148 1647 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00843 8185 3730 2335 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00842 2335 3735 2336 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00841 2334 2336 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00840 5182 7871 5184 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00839 8185 5184 5181 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00838 8185 7871 5185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00837 5183 5693 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00836 5184 5185 5183 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00835 8185 5180 5182 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00834 5181 5184 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00833 4359 5483 4358 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00832 4358 5654 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00831 4357 7353 4359 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00830 4552 7500 4357 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00829 6803 7345 6700 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00828 8185 7957 6805 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00827 6700 6805 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00826 8185 1807 962 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00825 845 962 961 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00824 8185 7314 845 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00823 963 961 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00822 8185 961 963 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00821 7582 7867 7856 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00820 8185 7856 7888 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00819 8185 7867 7857 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00818 7587 8058 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00817 7856 7857 7587 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00816 8185 7858 7582 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00815 7888 7856 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00814 7594 7867 7859 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00813 8185 7859 8186 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00812 8185 7867 7860 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00811 7595 8122 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00810 7859 7860 7595 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00809 8185 8119 7594 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00808 8186 7859 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00807 7589 7867 7590 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00806 8185 7590 7619 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00805 8185 7867 7593 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00804 7592 7591 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00803 7590 7593 7592 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00802 8185 7596 7589 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00801 7619 7590 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00800 8185 2006 2010 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00799 2010 2707 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00798 2011 2010 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00797 1242 1358 1241 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00796 1241 3819 1360 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00795 8185 1359 1242 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00794 1357 1360 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00793 2610 2614 2513 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00792 2513 3725 2610 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00791 8185 3315 2513 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00790 3038 3744 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00789 3100 3104 3038 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00788 3037 3102 3100 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00787 8185 3737 3037 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00786 3037 3098 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00785 8185 3556 2533 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00784 2646 2638 2530 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00783 2640 2648 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_00782 2530 2641 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00781 8185 3556 2641 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_00780 3567 2646 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_00779 2533 2642 2531 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00778 2531 2648 2646 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00777 2646 2640 2532 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00776 2532 3330 2533 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00775 6271 6974 6196 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00774 8185 7500 6272 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00773 6196 6272 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00772 7611 7867 7614 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00771 8185 7614 7630 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00770 8185 7867 7615 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00769 7613 7612 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00768 7614 7615 7613 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00767 8185 8137 7611 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00766 7630 7614 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00765 7609 7867 7865 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00764 8185 7865 8187 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00763 8185 7867 7866 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00762 7610 8139 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00761 7865 7866 7610 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00760 8185 8147 7609 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00759 8187 7865 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00758 3903 4574 3904 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00757 3904 7356 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00756 3902 6293 3903 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00755 3993 3994 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_00754 3994 6775 3902 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00753 2351 2827 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00752 2621 3307 2351 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00751 8185 2616 2621 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00750 8185 3556 2385 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00749 2387 2379 2381 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00748 2384 2648 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_00747 2381 2380 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00746 8185 3556 2380 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_00745 2845 2387 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_00744 2385 2382 2383 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00743 2383 2648 2387 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00742 2387 2384 2386 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00741 2386 3127 2385 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00740 3511 4885 3428 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00739 3428 5078 3511 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00738 8185 3765 3428 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00737 7236 7399 7237 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00736 7237 8176 7397 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00735 8185 7400 7236 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00734 7300 7397 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00733 8185 2202 1779 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00732 1657 1779 1777 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00731 8185 1780 1657 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00730 1778 1777 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00729 8185 1777 1778 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00728 7764 7766 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00727 8185 7787 7764 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00726 7764 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00725 8185 8045 7764 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00724 7765 7764 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00723 6207 7513 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00722 6288 6285 6207 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00721 6206 6286 6288 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00720 8185 6489 6206 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00719 6205 6349 6288 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00718 8185 6284 6205 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00717 7501 7754 7502 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00716 7502 7742 7501 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00715 8185 7500 7502 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00714 7741 7501 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00713 2373 4255 2374 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00712 2372 2371 2373 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00711 2374 3780 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00710 2631 2373 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00709 8185 2379 2372 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00708 2372 2840 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00707 2793 2795 3964 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00706 8185 3287 2793 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00705 2792 2794 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00704 3964 2791 2792 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00703 8185 2794 2795 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00702 2791 3287 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00701 6504 6506 6203 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00700 8185 7957 6282 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00699 6203 6282 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00698 8185 3723 2808 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00697 2808 2806 2807 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00696 2805 2807 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00695 8185 7026 1232 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00694 1232 6543 1349 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00693 2210 1349 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00692 4742 4734 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00691 5178 5664 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00690 6867 7957 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00689 4739 5863 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00688 6586 6870 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00687 8185 4075 3840 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00686 3840 3839 3843 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00685 3841 3843 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00684 799 2132 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00683 1292 1451 799 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00682 798 1929 1292 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00681 8185 1287 798 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00680 798 2595 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00679 6088 6087 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00678 6086 6083 6088 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00677 8185 6084 6086 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00676 6085 6086 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00675 6295 6821 6212 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00674 6212 6294 6295 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00673 8185 6297 6212 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00672 8185 4518 2097 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_00671 2097 2698 8185 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_00670 2236 2228 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00669 2097 5148 2228 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_00668 2228 2926 2097 8185 nmos_3p3 L=0.28U W=1.72U AS=0.4816P AD=0.4816P PS=4.01U PD=4.01U 
Mtr_00667 8185 3410 3034 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00666 3034 3182 3183 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00665 3261 3183 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00664 4722 4720 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00663 4731 4538 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00662 6142 6141 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00661 6358 6618 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00660 6381 6143 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00659 36 161 38 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00658 38 165 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00657 37 551 36 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00656 1114 158 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_00655 158 349 37 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00654 6063 7979 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00653 6062 6285 6063 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00652 6061 6286 6062 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00651 8185 6484 6061 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00650 6060 6292 6062 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00649 8185 6284 6060 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00648 7738 7802 7654 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00647 7654 7747 7738 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00646 8185 7737 7654 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00645 8185 8064 2788 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00644 2786 2788 2787 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00643 8185 5906 2786 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00642 3507 2787 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00641 8185 2787 3507 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00640 1783 7548 1659 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00639 1659 7559 1783 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00638 8185 1891 1659 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00637 1782 1783 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00636 2683 2682 2551 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00635 2552 4067 2683 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00634 2551 6796 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00633 7779 2683 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00632 8185 2898 2552 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00631 2552 2894 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00630 1598 6802 1599 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00629 1599 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00628 1596 6543 1598 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00627 1597 1595 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_00626 1595 5624 1596 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00625 3826 5453 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00624 8185 8159 3826 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00623 4281 6543 4282 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00622 4282 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00621 4279 5942 4281 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00620 4280 4278 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_00619 4278 7051 4279 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00618 1204 1297 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00617 3750 1298 1204 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00616 53 174 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00615 52 175 173 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00614 51 176 169 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00613 8185 4538 51 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00612 8185 3834 176 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00611 175 176 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00610 8185 177 174 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00609 173 176 53 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00608 170 173 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00607 8185 170 52 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00606 169 175 170 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00605 4538 169 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00604 8185 169 4538 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00603 7183 7348 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00602 7182 7350 7347 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00601 7181 7351 7344 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00600 8185 7345 7181 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00599 8185 8063 7351 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00598 7350 7351 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00597 8185 7349 7348 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00596 7347 7351 7183 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00595 7346 7347 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00594 8185 7346 7182 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00593 7344 7350 7346 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00592 7345 7344 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00591 8185 7344 7345 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00590 6042 6484 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00589 6260 6480 6042 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00588 8185 6481 6260 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00587 8185 7358 7464 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00586 7464 7359 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00585 8185 7357 7464 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00584 8185 3167 3168 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00583 3032 3168 3166 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00582 8185 3165 3032 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00581 3260 3166 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00580 8185 3166 3260 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00579 8185 7458 7507 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00578 7507 7514 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00577 7734 7507 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00576 408 509 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00575 407 510 507 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00574 406 511 506 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00573 8185 900 406 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00572 8185 1951 511 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00571 510 511 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00570 8185 899 509 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00569 507 511 408 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00568 505 507 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00567 8185 505 407 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00566 506 510 505 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00565 900 506 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00564 8185 506 900 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00563 7454 7725 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00562 7480 7724 7454 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00561 5835 5910 5758 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00560 5758 5911 5835 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00559 8185 5909 5758 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00558 7652 7733 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00557 7731 7742 7652 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00556 8185 7956 7731 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00555 7975 7731 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00554 6709 6830 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00553 6708 6833 6827 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00552 6707 6832 6824 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00551 8185 6823 6707 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00550 8185 8063 6832 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00549 6833 6832 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00548 8185 6829 6830 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00547 6827 6832 6709 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00546 6826 6827 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00545 8185 6826 6708 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00544 6824 6833 6826 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00543 6823 6824 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00542 8185 6824 6823 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00541 7987 7986 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00540 7983 7988 7984 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00539 7981 7989 7980 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00538 8185 7979 7981 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00537 8185 8063 7989 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00536 7988 7989 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00535 8185 7985 7986 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00534 7984 7989 7987 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00533 7982 7984 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00532 8185 7982 7983 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00531 7980 7988 7982 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00530 7979 7980 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00529 8185 7980 7979 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00528 8069 8067 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00527 8109 8068 8069 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00526 8185 7368 7471 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00525 7471 7369 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00524 8185 7367 7471 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00523 6640 6652 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00522 6639 6636 6640 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00521 1668 4575 1669 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00520 1669 2719 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00519 1813 4302 1668 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00518 5167 5169 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00517 5166 5168 5167 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00516 8185 6850 5166 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00515 5164 5166 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00514 1944 3542 1942 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00513 1942 2796 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00512 1943 3348 1944 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00511 2338 2346 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00510 2339 2610 2338 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00509 8185 2616 2339 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00508 2337 2339 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00507 6562 6564 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00506 6561 6565 6560 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00505 6557 6566 6558 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00504 8185 6567 6557 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00503 8185 8063 6566 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00502 6565 6566 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00501 8185 6563 6564 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00500 6560 6566 6562 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00499 6559 6560 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00498 8185 6559 6561 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00497 6558 6565 6559 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00496 6567 6558 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00495 8185 6558 6567 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00494 8185 4735 4352 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00493 4352 4744 4539 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00492 4447 4539 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00491 8185 6070 6072 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00490 6072 6071 6073 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00489 6332 6073 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00488 7217 7884 7218 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00487 7218 7398 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00486 7301 7883 7217 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00485 7115 7408 7113 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00484 7113 7881 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00483 7114 7883 7115 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00482 6534 6532 6533 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00481 6531 7550 6534 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00480 6533 6803 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00479 6530 6534 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00478 8185 7548 6531 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00477 6531 7559 8185 8185 nmos_3p3 L=0.28U W=2.88U AS=0.8064P AD=0.8064P PS=6.32U PD=6.32U 
Mtr_00476 2575 4575 2574 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00475 2574 2719 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00474 3404 2718 2575 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00473 2568 4575 2569 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00472 2569 2719 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00471 2925 4306 2568 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00470 8185 7330 7176 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00469 7176 7332 7331 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00468 7737 7331 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00467 2053 3566 2054 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00466 2054 3293 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00465 2152 3348 2053 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00464 3746 4512 3745 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00463 3745 4511 3747 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00462 8185 3744 3746 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00461 3743 3747 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00460 2869 3141 2870 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00459 8185 2870 2868 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00458 8185 3141 2872 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00457 2871 3348 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00456 2870 2872 2871 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00455 8185 3315 2869 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00454 2868 2870 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00453 4682 4684 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00452 4618 4620 4619 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00451 4616 4683 4680 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00450 8185 6549 4616 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00449 8185 8063 4683 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00448 4620 4683 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00447 8185 4681 4684 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00446 4619 4683 4682 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00445 4617 4619 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00444 8185 4617 4618 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00443 4680 4620 4617 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00442 6549 4680 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00441 8185 4680 6549 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00440 7504 7750 7505 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00439 7505 7747 7504 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00438 8185 7793 7505 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00437 7503 7504 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00436 4347 4529 4346 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00435 4346 4707 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00434 4345 4548 4347 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00433 5628 4527 4345 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00432 7150 7301 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00431 8185 7305 7150 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00430 7150 7147 7148 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00429 7148 7158 7150 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00428 7157 8187 7159 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00427 7159 7892 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00426 7158 7891 7157 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00425 7108 7114 7107 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00424 7107 7106 7108 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00423 8185 7104 7107 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00422 7621 8186 7620 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00421 7620 7619 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00420 7885 7869 7621 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00419 5263 7130 5261 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00418 5261 7887 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00417 5262 7149 5263 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00416 3796 4203 3795 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00415 3795 3794 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00414 4024 5908 3796 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00413 3292 4172 3294 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00412 3294 4173 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00411 3293 7528 3292 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00410 3911 5648 3910 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00409 3910 6797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00408 3909 6544 3911 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00407 4007 5603 3909 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00406 7213 7892 7214 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00405 7214 7398 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00404 7296 7869 7213 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00403 3800 7058 3799 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00402 3799 3797 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00401 3798 3801 3800 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00400 8048 5908 3798 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00399 2931 7356 2930 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00398 2930 4575 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00397 2929 4574 2931 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00396 3033 6293 2929 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00395 8061 8059 8060 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00394 8185 8064 8065 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00393 8060 8065 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00392 4328 4494 5092 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00391 8185 4497 4328 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00390 4329 4498 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00389 5092 4495 4329 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00388 8185 4498 4494 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00387 4495 4497 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00386 4514 5417 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00385 8185 7787 4514 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00384 4514 8048 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00383 8185 4429 4514 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00382 4428 4514 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00381 5247 6921 5248 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00380 5248 6172 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00379 5246 5868 5247 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00378 5245 7130 5246 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00377 4370 4573 4371 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00376 4371 4575 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00375 4369 4572 4370 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00374 4577 4574 4369 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00373 7232 7970 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00372 7263 7957 7232 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00371 4956 6090 4840 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00370 4840 6089 4956 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00369 8185 4955 4840 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00368 4677 5938 4679 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00367 4679 5108 4676 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00366 8185 5606 4677 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00365 4921 4676 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00364 5913 7787 5757 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00363 5757 5907 5913 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00362 8185 6801 5757 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00361 3410 3409 3411 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00360 3411 4779 3410 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00359 8185 3857 3411 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00358 8050 8055 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00357 8051 8064 8050 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00356 8185 4540 2915 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00355 2915 3379 2916 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00354 2918 2916 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00353 3312 3309 4914 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00352 8185 3310 3312 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00351 3314 3313 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00350 4914 3311 3314 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00349 8185 3313 3309 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00348 3311 3310 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00347 8185 8145 7868 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00346 7891 7868 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00345 8185 7868 7891 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00344 8185 7868 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00343 8144 7868 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00342 8185 8145 7864 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00341 7883 7864 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00340 8185 7864 7883 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00339 8185 7864 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00338 8144 7864 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00337 8185 8145 8146 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00336 8184 8146 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00335 8185 8146 8184 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00334 8185 8146 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00333 8144 8146 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00332 8185 8145 7870 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00331 7869 7870 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00330 8185 7870 7869 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00329 8185 7870 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00328 8144 7870 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00327 8185 5680 5681 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00326 8145 5681 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00325 8185 5681 8145 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00324 8185 5681 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00323 8144 5681 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00322 3408 4276 3407 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00321 3407 3405 3406 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00320 8185 3404 3408 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00319 3641 3406 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00318 2940 3857 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00317 3177 2943 2940 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00316 2939 4575 3177 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00315 8185 2937 2939 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00314 2939 2938 8185 8185 nmos_3p3 L=0.28U W=2.67U AS=0.7476P AD=0.7476P PS=5.9U PD=5.9U 
Mtr_00313 8185 1157 435 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00312 435 1372 564 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00311 565 564 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00310 1959 1956 1958 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00309 1958 1957 1959 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00308 8185 1962 1958 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00307 2167 1959 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00306 8185 969 573 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00305 5483 573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00304 8185 573 5483 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00303 8185 573 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00302 8144 573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00301 8185 969 970 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00300 5942 970 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00299 8185 970 5942 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00298 8185 970 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00297 8144 970 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00296 8185 579 578 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00295 969 578 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00294 8185 578 969 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00293 8185 578 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00292 8144 578 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00291 8185 384 382 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00290 5654 382 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00289 8185 382 5654 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00288 8185 382 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00287 8144 382 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00286 8185 384 383 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00285 5447 383 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00284 8185 383 5447 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00283 8185 383 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00282 8144 383 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00281 8185 386 385 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00280 384 385 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00279 8185 385 384 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00278 8185 385 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00277 8144 385 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00276 8185 6312 6313 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00275 7352 6313 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00274 8185 6313 7352 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00273 8185 6313 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00272 8144 6313 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00271 8185 6312 6306 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00270 7041 6306 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00269 8185 6306 7041 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00268 8185 6306 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00267 8144 6306 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00266 8185 5916 5915 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00265 6312 5915 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00264 8185 5915 6312 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00263 8185 5915 8144 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00262 8144 5915 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00261 5442 5444 5314 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00260 5314 5633 5442 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00259 8185 7068 5314 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00258 5440 5442 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00257 3468 3801 3469 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00256 3469 7058 3605 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00255 8185 5908 3468 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00254 5633 3605 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00253 1590 1377 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00252 8185 1375 1590 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00251 4879 5037 4880 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00250 4880 5509 5039 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00249 8185 5038 4879 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00248 5036 5039 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00247 1577 2022 1578 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00246 1578 1583 1579 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00245 8185 1576 1577 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00244 3156 1579 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00243 4194 4192 4195 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00242 4195 4193 4196 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00241 8185 4438 4194 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00240 4191 4196 8185 8185 nmos_3p3 L=0.28U W=2.98U AS=0.8344P AD=0.8344P PS=6.53U PD=6.53U 
Mtr_00239 2883 6076 2882 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00238 8185 8064 2884 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00237 2882 2884 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00236 4661 4659 4662 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00235 8185 4658 4661 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00234 4664 4663 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00233 4662 4660 4664 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00232 8185 4663 4659 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00231 4660 4658 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00230 840 4068 841 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00229 841 6311 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00228 839 4572 840 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00227 1375 959 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_00226 959 3857 839 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00225 814 932 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00224 813 933 931 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00223 812 934 927 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00222 8185 1113 812 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00221 8185 3834 934 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00220 933 934 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00219 8185 935 932 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00218 931 934 814 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00217 929 931 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00216 8185 929 813 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00215 927 933 929 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00214 1113 927 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00213 8185 927 1113 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00212 8185 6127 5854 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00211 5854 6145 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00210 8185 6618 5854 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00209 7790 7791 7664 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00208 7664 7788 7790 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00207 8185 8040 7664 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00206 7789 7790 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00205 1187 4068 1189 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00204 1189 4295 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00203 1188 5648 1187 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00202 1390 1186 8185 8185 nmos_3p3 L=0.28U W=2.56U AS=0.7168P AD=0.7168P PS=5.69U PD=5.69U 
Mtr_00201 1186 4067 1188 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00200 1619 1617 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00199 8185 1618 1619 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00198 8185 3650 3268 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00197 3268 3664 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00196 8185 3267 3268 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00195 4753 4754 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00194 4632 4634 4633 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00193 4630 4755 4752 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00192 8185 4760 4630 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00191 8185 5864 4755 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00190 4634 4755 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00189 8185 4759 4754 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00188 4633 4755 4753 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00187 4631 4633 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00186 8185 4631 4632 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00185 4752 4634 4631 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00184 4760 4752 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00183 8185 4752 4760 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00182 4735 4734 4736 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00181 4736 6363 4735 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00180 8185 6359 4736 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00179 4239 4449 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00178 4244 4448 4239 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00177 5800 7633 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00176 6156 6396 5800 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00175 5351 7633 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00174 6158 6652 5351 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00173 7673 7820 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00172 7672 7822 7818 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00171 7671 7823 7814 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00170 8185 8071 7671 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00169 8185 7821 7823 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00168 7822 7823 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00167 8185 8070 7820 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00166 7818 7823 7673 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00165 7817 7818 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00164 8185 7817 7672 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00163 7814 7822 7817 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00162 8071 7814 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00161 8185 7814 8071 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00160 7523 7797 7524 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00159 7524 7798 7523 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00158 8185 8139 7524 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00157 5159 7352 5158 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00156 5158 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00155 5160 5435 5159 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00154 4397 4749 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00153 4448 4955 4397 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00152 6034 8179 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00151 6615 7872 6034 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00150 438 6609 439 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00149 439 1565 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00148 5148 4306 438 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00147 1259 6802 1258 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00146 1258 1565 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00145 4518 4306 1259 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00144 2957 2712 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00143 8185 2942 2957 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00142 2957 2932 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00141 8185 2710 2957 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00140 341 3622 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00139 342 1150 341 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00138 39 365 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00137 159 166 39 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00136 3007 3780 3147 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00135 8185 3147 3315 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00134 8185 3780 3070 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00133 3008 3353 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00132 3147 3070 3008 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00131 8185 3602 3007 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00130 3315 3147 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00129 3360 3780 3359 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00128 8185 3359 4510 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00127 8185 3780 3363 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00126 3362 3361 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00125 3359 3363 3362 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00124 8185 5180 3360 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00123 4510 3359 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00122 3351 3780 3350 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00121 8185 3350 3348 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00120 8185 3780 3355 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00119 3354 3353 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00118 3350 3355 3354 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00117 8185 4030 3351 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00116 3348 3350 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00115 5564 7041 5565 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00114 5565 7361 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00113 5562 5563 5564 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00112 5347 5498 8185 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00111 5495 5706 5347 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00110 1248 6609 1249 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00109 1249 4068 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00108 1543 6796 1248 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00107 8185 1466 1468 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00106 1468 5099 1469 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00105 1467 1469 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00104 8185 2798 2507 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00103 2507 3553 2600 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00102 2599 2600 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00101 8185 3556 3443 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00100 3549 3757 3441 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00099 3547 3562 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_00098 3441 3545 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00097 8185 3556 3545 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_00096 3986 3549 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_00095 3443 3546 3442 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00094 3442 3562 3549 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00093 3549 3547 3444 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00092 3444 4426 3443 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00091 8185 3556 3448 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00090 3563 3995 3446 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00089 3560 3562 8185 8185 nmos_3p3 L=0.28U W=0.78U AS=0.2184P AD=0.2184P PS=2.12U PD=2.12U 
Mtr_00088 3446 3558 8185 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00087 8185 3556 3558 8185 nmos_3p3 L=0.28U W=0.57U AS=0.1596P AD=0.1596P PS=1.7U PD=1.7U 
Mtr_00086 4141 3563 8185 8185 nmos_3p3 L=0.28U W=2.77U AS=0.7756P AD=0.7756P PS=6.11U PD=6.11U 
Mtr_00085 3448 3559 3447 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00084 3447 3562 3563 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00083 3563 3560 3449 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00082 3449 3754 3448 8185 nmos_3p3 L=0.28U W=1.2U AS=0.336P AD=0.336P PS=2.96U PD=2.96U 
Mtr_00081 7994 7996 8185 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00080 7993 7997 7995 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00079 7990 7998 7991 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00078 8185 8000 7990 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00077 8185 8063 7998 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00076 7997 7998 8185 8185 nmos_3p3 L=0.28U W=1.41U AS=0.3948P AD=0.3948P PS=3.38U PD=3.38U 
Mtr_00075 8185 7999 7996 8185 nmos_3p3 L=0.28U W=1.83U AS=0.5124P AD=0.5124P PS=4.22U PD=4.22U 
Mtr_00074 7995 7998 7994 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00073 7992 7995 8185 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00072 8185 7992 7993 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00071 7991 7997 7992 8185 nmos_3p3 L=0.28U W=0.99U AS=0.2772P AD=0.2772P PS=2.54U PD=2.54U 
Mtr_00070 8000 7991 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00069 8185 7991 8000 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00068 6784 5417 5299 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00067 5299 5432 6784 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00066 8185 5416 5299 8185 nmos_3p3 L=0.28U W=2.04U AS=0.5712P AD=0.5712P PS=4.64U PD=4.64U 
Mtr_00065 8185 4518 2093 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00064 2093 2227 2219 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00063 2437 2219 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00062 7401 8180 7219 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00061 7219 7639 7401 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00060 8185 7633 7219 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00059 7302 7401 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00058 6572 6867 6573 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00057 8185 6573 6843 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00056 8185 6867 6575 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00055 6574 6663 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00054 6573 6575 6574 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00053 8185 6838 6572 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00052 6843 6573 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00051 6719 6867 6866 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00050 8185 6866 6863 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00049 8185 6867 6869 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00048 6720 7283 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00047 6866 6869 6720 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00046 8185 6864 6719 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00045 6863 6866 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00044 6603 6867 6605 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00043 8185 6605 6600 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00042 8185 6867 6606 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00041 6604 6632 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00040 6605 6606 6604 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00039 8185 6602 6603 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00038 6600 6605 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00037 54 4538 179 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00036 8185 179 177 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00035 8185 4538 181 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00034 55 187 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00033 179 181 55 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00032 8185 4540 54 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00031 177 179 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00030 6731 7867 6902 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00029 8185 6902 6900 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00028 8185 7867 6904 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00027 6732 6988 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00026 6902 6904 6732 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00025 8185 7119 6731 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00024 6900 6902 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00023 7208 7867 7387 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00022 8185 7387 7893 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00021 8185 7867 7292 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00020 7209 7777 8185 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00019 7387 7292 7209 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00018 8185 7604 7208 8185 nmos_3p3 L=0.28U W=0.88U AS=0.2464P AD=0.2464P PS=2.33U PD=2.33U 
Mtr_00017 7893 7387 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00016 1982 5648 1983 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00015 1983 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00014 4517 7051 1982 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00013 829 5483 830 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00012 830 4310 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00011 5147 7051 829 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00010 8185 7343 6688 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00009 6688 6794 6791 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00008 7007 6791 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00007 1933 2152 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00006 1932 2608 1933 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00005 8185 2616 1932 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00004 2518 2827 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00003 2617 3307 2518 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00002 8185 2616 2617 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
Mtr_00001 2816 2617 8185 8185 nmos_3p3 L=0.28U W=1.93U AS=0.5404P AD=0.5404P PS=4.43U PD=4.43U 
.ends arlet6502_cts_r

