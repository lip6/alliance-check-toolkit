* Spice description of ao22_x2
* Spice driver version 1456475931
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:34

* INTERF i0 i1 i2 q vdd vss 


.subckt ao22_x2 7 6 3 4 2 5 
* NET 2 = vdd
* NET 3 = i2
* NET 4 = q
* NET 5 = vss
* NET 6 = i1
* NET 7 = i0
Mtr_00008 4 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00007 2 3 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00006 1 7 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00005 8 6 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00004 4 8 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 5 3 9 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 9 6 8 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 8 7 9 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C8 2 5 1.97889e-15
C7 3 5 2.3779e-15
C6 4 5 2.22185e-15
C5 5 5 1.87591e-15
C4 6 5 1.68468e-15
C3 7 5 1.39432e-15
C2 8 5 2.01414e-15
C1 9 5 4.9821e-16
.ends ao22_x2

