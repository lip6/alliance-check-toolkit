* pnp_t
.param
+ dkispp=9.2840e-01 dkbfpp=9.5154e-01 dknfpp=1.000
+ dkispp5x=1.0046e+00 dkbfpp5x=1.1288e+00 dknfpp5x=1.0009e+00 dkisepp5x=0.745
