* Spice description of oa2a2a2a24_x4
* Spice driver version 1867521819
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:32

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss 


.subckt oa2a2a2a24_x4 5 4 8 9 11 12 13 16 6 1 18 
* NET 1 = vdd
* NET 4 = i1
* NET 5 = i0
* NET 6 = q
* NET 8 = i2
* NET 9 = i3
* NET 11 = i4
* NET 12 = i5
* NET 13 = i6
* NET 16 = i7
* NET 18 = vss
Mtr_00020 1 15 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00019 6 15 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00018 1 5 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00017 2 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00016 3 8 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 2 9 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 3 11 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 3 12 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 3 13 15 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 15 16 3 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 7 4 15 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4488P AD=0.4488P PS=4.22U PD=4.22U 
Mtr_00009 6 15 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4488P AD=0.4488P PS=4.22U PD=4.22U 
Mtr_00008 18 5 7 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4488P AD=0.4488P PS=4.22U PD=4.22U 
Mtr_00007 18 15 6 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4488P AD=0.4488P PS=4.22U PD=4.22U 
Mtr_00006 18 8 10 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 10 9 15 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 15 11 14 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 14 12 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 15 13 17 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 17 16 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C18 1 18 4.65318e-15
C17 2 18 7.56633e-16
C16 3 18 2.39396e-15
C15 4 18 1.40338e-15
C14 5 18 1.38512e-15
C13 6 18 1.80209e-15
C11 8 18 1.43912e-15
C10 9 18 1.42999e-15
C8 11 18 1.43912e-15
C7 12 18 1.43912e-15
C6 13 18 1.46243e-15
C4 15 18 3.63534e-15
C3 16 18 1.74315e-15
C1 18 18 3.84163e-15
.ends oa2a2a2a24_x4

