* Spice description of xr2_x1
* Spice driver version 101932827
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:44

* INTERF i0 i1 q vdd vss 


.subckt xr2_x1 7 3 6 1 9 
* NET 1 = vdd
* NET 3 = i1
* NET 6 = q
* NET 7 = i0
* NET 9 = vss
Mtr_00012 2 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00011 1 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 1 8 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 6 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 1 7 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 7 8 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00006 4 8 6 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 9 2 4 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 2 3 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 5 7 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 6 3 5 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 9 7 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C9 1 9 3.34343e-15
C8 2 9 2.23e-15
C7 3 9 3.32219e-15
C4 6 9 2.08504e-15
C3 7 9 2.63951e-15
C2 8 9 1.853e-15
C1 9 9 2.20432e-15
.ends xr2_x1

