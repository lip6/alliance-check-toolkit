* tie
.subckt tie vdd vss

.ends tie
