* Spice description of noa2a22_x1
* Spice driver version -381931749
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:07

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt noa2a22_x1 8 7 4 3 6 1 10 
* NET 1 = vdd
* NET 3 = i3
* NET 4 = i2
* NET 6 = nq
* NET 7 = i1
* NET 8 = i0
* NET 10 = vss
Mtr_00008 2 4 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 3 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00006 2 7 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 6 8 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 5 3 6 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 6 7 9 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 10 4 5 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 9 8 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C10 1 10 1.66309e-15
C9 2 10 8.0812e-16
C8 3 10 2.10592e-15
C7 4 10 2.14834e-15
C5 6 10 2.03943e-15
C4 7 10 1.70741e-15
C3 8 10 1.70741e-15
C1 10 10 1.71458e-15
.ends noa2a22_x1

