* inv_x2
* inv_x2
.subckt inv_x2 vdd vss i nq
Mnmos[0] vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[0] vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
Mnmos[1] nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.735um
Mpmos[1] nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.295um
.ends inv_x2
