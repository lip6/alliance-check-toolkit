* Spice description of inv_x1
* Spice driver version 2051432219
* Date ( dd/mm/yyyy hh:mm:ss ):  9/07/2024 at 14:35:08

* INTERF i nq vdd vss 


.subckt inv_x1 2 4 1 3 
* NET 1 = vdd
* NET 2 = i
* NET 3 = vss
* NET 4 = nq
Mtr_00002 4 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_00001 4 2 3 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
.ends inv_x1

