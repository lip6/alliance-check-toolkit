-- no model for inv_x0
