* pnp_s
.param
+ dkispp=7.0967e-01 dkbfpp=4.9061e-01 dknfpp=1.000
+ dkispp5x=7.8658e-01 dkbfpp5x=4.6158e-01 dknfpp5x=1.0009e+00 dkisepp5x=0.745
