* rc_model
.model sky130_fd_pr__res_generic_nd r tc1r={tc1rsn} tc2r={tc2rsn} rsh={rdn} dw={-tol_nfom/2-nfom_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_pd r tc1r={tc1rsp} tc2r={tc2rsp} rsh={rdp} dw={-tol_pfom/2-pfom_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_nd__hv r tc1r={tc1rsn_h} tc2r={tc2rsn_h} rsh={rdn_hv} dw={-tol_nfom/2-nfom_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_pd__hv r tc1r={tc1rsp_h} tc2r={tc2rsp_h} rsh={rdp_hv} dw={-tol_pfom/2-pfom_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_po r tc1r=tc1rsgpu tc2r=tc2rsgpu rsh=rp1 dw={-tol_poly/2-poly_dw/2} tnom=30
.model sky130_fd_pr__res_generic_nw r tc1r={tc1rsnw} tc2r={tc2rsnw} rsh={rnw} dw={-tol_nw/2} tnom=30.0
.model sky130_fd_pr__res_generic_l1 r tc1r={tc1rl1} tc2r={tc2rl1} rsh={rl1} dw={-tol_li/2-li_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_m1 r tc1r={tc1rm1} tc2r={tc2rm1} rsh={rm1} dw={-tol_m1/2-m1_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_m2 r tc1r={tc1rm2} tc2r={tc2rm2} rsh={rm2} dw={-tol_m2/2-m2_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_m3 r tc1r={tc1rm3} tc2r={tc2rm3} rsh={rm3} dw={-tol_m3/2-m3_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_m4 r tc1r={tc1rm4} tc2r={tc2rm4} rsh={rm4} dw={-tol_m4/2-m4_dw/2} tnom=30.0
.model sky130_fd_pr__res_generic_m5 r tc1r={tc1rm5} tc2r={tc2rm5} rsh={rm5} dw={-tol_m5/2-m5_dw/2} tnom=30.0
