*
* sky130_fd_sc_hd__inv_1_chain.spi
* 

* sky130_fd_sc_hd__inv_1
*.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y

.INCLUDE sky130_fd_sc_hd__inv_1.spice

.subckt sky130_fd_sc_hd__inv_1_chain in out vdd gnd
Xa in gnd gnd vdd vdd n1   sky130_fd_sc_hd__inv_1
Xb n1 gnd gnd vdd vdd n2   sky130_fd_sc_hd__inv_1
Xc n2 gnd gnd vdd vdd n3   sky130_fd_sc_hd__inv_1
Xd n3 gnd gnd vdd vdd n4   sky130_fd_sc_hd__inv_1
Xe n4 gnd gnd vdd vdd n5   sky130_fd_sc_hd__inv_1
Xf n5 gnd gnd vdd vdd n6   sky130_fd_sc_hd__inv_1
Xg n6 gnd gnd vdd vdd n7   sky130_fd_sc_hd__inv_1
Xh n7 gnd gnd vdd vdd n8   sky130_fd_sc_hd__inv_1
Xi n8 gnd gnd vdd vdd n9   sky130_fd_sc_hd__inv_1
Xj n9 gnd gnd vdd vdd out  sky130_fd_sc_hd__inv_1
.ends sky130_fd_sc_hd__inv_1_chain


