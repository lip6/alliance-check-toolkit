* Filler400
.subckt Filler400 vss vdd iovss iovdd

.ends Filler400
