-- no model for inv_x4
