* Spice description of inv_x2
* Spice driver version -114258149
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:41

* INTERF i nq vdd vss 


.subckt inv_x2 2 4 1 3 
* NET 1 = vdd
* NET 2 = i
* NET 3 = vss
* NET 4 = nq
Mtr_00002 4 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00001 4 2 3 3 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
C4 1 3 1.27468e-15
C3 2 3 1.65586e-15
C2 3 3 1.19279e-15
C1 4 3 2.23361e-15
.ends inv_x2

