../rtl/snx.vhdl