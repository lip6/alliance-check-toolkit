* Spice description of noa2a2a2a24_x1
* Spice driver version -271180005
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:11

* INTERF i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss 


.subckt noa2a2a2a24_x1 6 5 8 9 11 12 13 16 15 2 18 
* NET 2 = vdd
* NET 5 = i1
* NET 6 = i0
* NET 8 = i2
* NET 9 = i3
* NET 11 = i4
* NET 12 = i5
* NET 13 = i6
* NET 15 = nq
* NET 16 = i7
* NET 18 = vss
Mtr_00016 1 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00015 2 6 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00014 1 9 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 3 8 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 3 11 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 4 12 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 4 13 15 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 15 16 4 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 7 5 15 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00007 18 6 7 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00006 18 8 10 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00005 10 9 15 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00004 15 11 14 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00003 14 12 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00002 15 13 17 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
Mtr_00001 17 16 18 18 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.53U AS=0.3672P AD=0.3672P PS=3.54U PD=3.54U 
C18 1 18 8.93446e-16
C17 2 18 3.10802e-15
C16 3 18 1.01162e-15
C15 4 18 1.35193e-15
C14 5 18 1.38512e-15
C13 6 18 1.68915e-15
C11 8 18 1.43826e-15
C10 9 18 1.42913e-15
C8 11 18 1.43344e-15
C7 12 18 1.45169e-15
C6 13 18 1.4431e-15
C4 15 18 2.85099e-15
C3 16 18 1.77505e-15
C1 18 18 3.19392e-15
.ends noa2a2a2a24_x1

