*
* 

*****************

.TEMP 25

******************
* BSIM4 transistor model parameters for ngspice
*.lib /users/soft/analogdesign/scalable/techno/sky130_models_20220217/C4M.Sky130_all_lib.spice logic_tt 

*******************************
*Simulation conditions

Vground evss 0 0
Vsupply evdd 0 DC 1.8
*gfoncd evdd 0 evdd 0 1.0e-15

******************
* circuit model
* include circuit netlist
.include mac_cts_r.spi
*****************

*****************
* Circuit Instantiation
*.subckt inv_x2 vdd vss i nq

Xc evss evdd 23 32 33 34 35 36 37 38 39 93 95 96 97 98 99 100 101 102 mac_cts_r
.end

