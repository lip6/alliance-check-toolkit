-- no model for tie
