* Spice description of no4_x4
* Spice driver version -2025787621
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:04

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt no4_x4 8 10 7 9 6 3 12 
* NET 3 = vdd
* NET 6 = nq
* NET 7 = i2
* NET 8 = i0
* NET 9 = i3
* NET 10 = i1
* NET 12 = vss
Mtr_00014 5 11 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.78U AS=0.4272P AD=0.4272P PS=4.05U PD=4.05U 
Mtr_00013 3 5 6 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.4U AS=0.816P AD=0.816P PS=7.28U PD=7.28U 
Mtr_00012 6 5 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.4U AS=0.816P AD=0.816P PS=7.28U PD=7.28U 
Mtr_00011 3 9 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.4U AS=0.816P AD=0.816P PS=7.28U PD=7.28U 
Mtr_00010 1 7 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.4U AS=0.816P AD=0.816P PS=7.28U PD=7.28U 
Mtr_00009 2 8 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.4U AS=0.816P AD=0.816P PS=7.28U PD=7.28U 
Mtr_00008 4 10 11 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.4U AS=0.816P AD=0.816P PS=7.28U PD=7.28U 
Mtr_00007 11 10 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00006 11 7 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00005 12 9 11 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00004 12 8 11 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 6 5 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00002 12 5 6 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00001 5 11 12 12 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C10 3 12 3.35605e-15
C8 5 12 1.95907e-15
C7 6 12 1.99971e-15
C6 7 12 2.04794e-15
C5 8 12 2.0662e-15
C4 9 12 2.08445e-15
C3 10 12 2.02056e-15
C2 11 12 3.3497e-15
C1 12 12 2.85558e-15
.ends no4_x4

