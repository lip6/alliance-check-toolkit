* Spice description of oa2a22_x2
* Spice driver version -1081839845
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:27

* INTERF i0 i1 i2 i3 q vdd vss 


.subckt oa2a22_x2 9 8 5 4 3 2 11 
* NET 2 = vdd
* NET 3 = q
* NET 4 = i3
* NET 5 = i2
* NET 8 = i1
* NET 9 = i0
* NET 11 = vss
Mtr_00010 3 6 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 6 9 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 1 8 6 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 2 5 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 1 4 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 11 4 7 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00004 7 5 6 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00003 6 8 10 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 3 6 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 10 9 11 11 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C11 1 11 8.84127e-16
C10 2 11 2.7287e-15
C9 3 11 2.15173e-15
C8 4 11 1.88082e-15
C7 5 11 1.83894e-15
C6 6 11 2.63396e-15
C4 8 11 1.81961e-15
C3 9 11 1.51558e-15
C1 11 11 2.9322e-15
.ends oa2a22_x2

