* Spice description of oa3ao322_x2
* Spice driver version 81383195
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:35

* INTERF i0 i1 i2 i3 i4 i5 i6 q vdd vss 


.subckt oa3ao322_x2 12 11 10 7 5 6 8 16 4 17 
* NET 4 = vdd
* NET 5 = i4
* NET 6 = i5
* NET 7 = i3
* NET 8 = i6
* NET 10 = i2
* NET 11 = i1
* NET 12 = i0
* NET 16 = q
* NET 17 = vss
Mtr_00016 3 7 15 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00015 1 5 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00014 15 8 2 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00013 2 12 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00012 4 11 2 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00011 2 10 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00010 4 15 16 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 2 6 1 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00008 17 7 9 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00007 9 8 15 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.78U AS=0.4272P AD=0.4272P PS=4.05U PD=4.05U 
Mtr_00006 15 10 14 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00005 14 11 13 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00004 17 15 16 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.12U AS=0.5088P AD=0.5088P PS=4.73U PD=4.73U 
Mtr_00003 13 12 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.36U AS=0.3264P AD=0.3264P PS=3.2U PD=3.2U 
Mtr_00002 9 5 17 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
Mtr_00001 17 6 9 17 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.44U AS=0.3456P AD=0.3456P PS=3.37U PD=3.37U 
C16 2 17 1.26416e-15
C14 4 17 3.19392e-15
C13 5 17 1.69828e-15
C12 6 17 1.72566e-15
C11 7 17 1.68915e-15
C10 8 17 1.42163e-15
C9 9 17 6.56106e-16
C8 10 17 1.376e-15
C7 11 17 1.68002e-15
C6 12 17 1.69828e-15
C3 15 17 2.39102e-15
C2 16 17 2.15173e-15
C1 17 17 3.28512e-15
.ends oa3ao322_x2

