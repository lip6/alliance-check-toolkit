* Filler10000
.subckt Filler10000 vss vdd iovss iovdd

.ends Filler10000
