-- no model for buf_x1
