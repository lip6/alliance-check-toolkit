* Spice description of oa22_x2
* Spice driver version 1536663323
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:26

* INTERF i0 i1 i2 q vdd vss 


.subckt oa22_x2 7 6 3 4 2 9 
* NET 2 = vdd
* NET 3 = i2
* NET 4 = q
* NET 6 = i1
* NET 7 = i0
* NET 9 = vss
Mtr_00008 4 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 1 6 5 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 2 3 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00005 5 7 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00004 4 5 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 9 3 5 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 5 6 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 8 7 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C9 1 9 7.47315e-16
C8 2 9 1.66309e-15
C7 3 9 2.34743e-15
C6 4 9 2.15173e-15
C5 5 9 1.61286e-15
C4 6 9 1.70287e-15
C3 7 9 1.88995e-15
C1 9 9 1.71458e-15
.ends oa22_x2

