* Spice description of no3_x1
* Spice driver version 561471259
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:02

* INTERF i0 i1 i2 nq vdd vss 


.subckt no3_x1 5 6 4 8 2 7 
* NET 2 = vdd
* NET 4 = i2
* NET 5 = i0
* NET 6 = i1
* NET 7 = vss
* NET 8 = nq
Mtr_00006 2 4 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 1 5 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 3 6 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 7 4 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 8 5 7 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 7 6 8 7 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C7 2 7 1.41822e-15
C5 4 7 2.36378e-15
C4 5 7 1.75572e-15
C3 6 7 1.76538e-15
C2 7 7 1.57612e-15
C1 8 7 2.74971e-15
.ends no3_x1

