-- no model for or4_x1
