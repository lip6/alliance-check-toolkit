* Spice description of one_x0
* Spice driver version -2088358117
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:39

* INTERF q vdd vss 


.subckt one_x0 2 1 3 
* NET 1 = vdd
* NET 2 = q
* NET 3 = vss
Mtr_00001 2 3 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C3 1 3 1.43601e-15
C2 2 3 2.04875e-15
C1 3 3 1.6988e-15
.ends one_x0

