* IOPadVss
.subckt IOPadVss vss vdd iovss iovdd
Xpad vss Pad_15800W12000H
Xnclamp iovss iovdd vss Clamp_N32N0D
Xpclamp iovss iovdd vss Clamp_P32N0D
Xbulkconn vdd vss iovdd iovss BulkConn_18000WUp
.ends IOPadVss
