-- no model for mux2_x1
