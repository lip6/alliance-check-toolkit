-- no model for tie_poly
