* a2_x2
* a2_x2
.subckt a2_x2 vss q vdd i0 i1
Mn_net0_1 vss _net0 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net0_1 vdd _net0 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i0_1 _net0 i0 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i0_1 vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i1_1 _net0 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i1_1 _net1 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
.ends a2_x2
