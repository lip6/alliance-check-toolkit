* Spice description of nao2o22_x4
* Spice driver version 403164955
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:56

* INTERF i0 i1 i2 i3 nq vdd vss 


.subckt nao2o22_x4 10 7 6 8 4 3 9 
* NET 3 = vdd
* NET 4 = nq
* NET 6 = i2
* NET 7 = i1
* NET 8 = i3
* NET 9 = vss
* NET 10 = i0
Mtr_00014 4 5 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 3 5 4 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 1 8 11 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00011 2 10 3 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00010 3 6 1 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00009 11 7 2 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00008 3 11 5 3 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 4 5 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00006 9 5 4 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00005 12 6 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00004 12 7 11 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00003 11 10 12 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
Mtr_00002 9 11 5 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 9 8 12 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.19U AS=0.2856P AD=0.2856P PS=2.86U PD=2.86U 
C10 3 9 3.97601e-15
C9 4 9 2.15173e-15
C8 5 9 1.9814e-15
C7 6 9 1.84753e-15
C6 7 9 1.82874e-15
C5 8 9 1.85666e-15
C4 9 9 3.42782e-15
C3 10 9 1.79868e-15
C2 11 9 2.80086e-15
C1 12 9 8.68926e-16
.ends nao2o22_x4

