* Spice description of m65_cts_r_ext
* Spice driver version 492387240
* Date ( dd/mm/yyyy hh:mm:ss ): 10/07/2024 at 15:08:09

* INTERF adrs[0] adrs[1] adrs[2] adrs[3] adrs[4] adrs[5] adrs[6] adrs[7] 
* INTERF adrs[8] adrs[9] adrs[10] adrs[11] adrs[12] adrs[13] adrs[14] 
* INTERF adrs[15] data[0] data[1] data[2] data[3] data[4] data[5] data[6] 
* INTERF data[7] datao[0] datao[1] datao[2] datao[3] datao[4] datao[5] 
* INTERF datao[6] datao[7] debug[0] debug[1] debug[2] debug[3] debug[4] 
* INTERF debug[5] debug[6] debug[7] debug[8] debug[9] debug[10] debug[11] 
* INTERF debug[12] debug[13] debug[14] debug[15] irq m_clock nmi p_reset rd 
* INTERF rdy start sync vdd vss wt 


.subckt m65_cts_r_ext 5536 5523 6187 5969 5454 5746 5160 5833 4642 4975 5350 4959 5045 6539 7511 7495 5043 5055 5274 5216 4834 5137 4979 5138 5267 5812 7123 6762 6476 5991 5256 5540 7494 7493 7489 7481 7480 7475 7466 7464 7462 7454 7453 7452 7335 6965 6676 6628 4938 3717 6410 1412 1841 2754 1115 5623 7451 7514 6409 
* NET 11 = subckt_1662_sff1_x4.sff_s
* NET 13 = subckt_1662_sff1_x4.sff_m
* NET 17 = subckt_1662_sff1_x4.ckr
* NET 18 = subckt_1662_sff1_x4.nckr
* NET 33 = subckt_1574_sff1_x4.sff_s
* NET 36 = subckt_1574_sff1_x4.sff_m
* NET 38 = subckt_1574_sff1_x4.ckr
* NET 40 = subckt_1574_sff1_x4.nckr
* NET 41 = abc_8306_auto_rtlil_cc_2608_muxgate_8073
* NET 66 = subckt_1654_sff1_x4.sff_s
* NET 69 = subckt_1654_sff1_x4.sff_m
* NET 73 = subckt_1654_sff1_x4.ckr
* NET 74 = subckt_1654_sff1_x4.nckr
* NET 78 = abc_8306_new_n862
* NET 84 = subckt_1615_sff1_x4.sff_s
* NET 87 = subckt_1615_sff1_x4.sff_m
* NET 91 = subckt_1615_sff1_x4.ckr
* NET 92 = subckt_1615_sff1_x4.nckr
* NET 93 = subckt_1576_sff1_x4.sff_s
* NET 96 = subckt_1576_sff1_x4.sff_m
* NET 100 = subckt_1576_sff1_x4.ckr
* NET 101 = subckt_1576_sff1_x4.nckr
* NET 102 = subckt_1579_sff1_x4.sff_s
* NET 105 = subckt_1579_sff1_x4.sff_m
* NET 109 = subckt_1579_sff1_x4.ckr
* NET 110 = subckt_1579_sff1_x4.nckr
* NET 121 = subckt_1653_sff1_x4.sff_m
* NET 124 = subckt_1653_sff1_x4.ckr
* NET 125 = subckt_1653_sff1_x4.nckr
* NET 126 = abc_8306_new_n864
* NET 130 = abc_8306_auto_rtlil_cc_2608_muxgate_8077
* NET 132 = abc_8306_auto_rtlil_cc_2608_muxgate_8083
* NET 141 = subckt_1653_sff1_x4.sff_s
* NET 162 = abc_8306_new_n1295
* NET 181 = abc_8306_new_n825
* NET 186 = abc_8306_new_n767
* NET 190 = ex_st[2]
* NET 191 = ex_st_bit2_hfns_2
* NET 193 = abc_8306_new_n1299
* NET 195 = abc_8306_new_n444
* NET 225 = abc_8306_new_n776
* NET 230 = subckt_1578_sff1_x4.sff_s
* NET 233 = abc_8306_auto_rtlil_cc_2608_muxgate_8081
* NET 235 = subckt_1578_sff1_x4.sff_m
* NET 236 = subckt_1578_sff1_x4.ckr
* NET 238 = subckt_1578_sff1_x4.nckr
* NET 239 = abc_8306_new_n1305
* NET 242 = abc_8306_new_n443
* NET 262 = abc_8306_new_n1025
* NET 266 = abc_8306_new_n1033
* NET 272 = abc_8306_new_n802
* NET 275 = abc_8306_new_n851
* NET 276 = abc_8306_new_n863
* NET 280 = abc_8306_new_n871
* NET 281 = abc_8306_new_n768
* NET 283 = abc_8306_new_n784
* NET 286 = op[5]
* NET 290 = subckt_1573_sff1r_x4.sff_s
* NET 294 = subckt_1573_sff1r_x4.sff_m
* NET 295 = abc_8306_auto_rtlil_cc_2608_muxgate_8071
* NET 297 = subckt_1573_sff1r_x4.ckr
* NET 298 = subckt_1573_sff1r_x4.nckr
* NET 310 = spare_buffer_338.q
* NET 312 = abc_8306_new_n1104
* NET 316 = spare_buffer_334.q
* NET 320 = spare_buffer_322.q
* NET 325 = abc_8306_new_n773
* NET 326 = spare_buffer_318.q
* NET 329 = spare_buffer_258.q
* NET 331 = op_bit6_hfns_2
* NET 333 = spare_buffer_254.q
* NET 335 = spare_buffer_242.q
* NET 338 = abc_8306_new_n1297
* NET 340 = abc_8306_new_n337
* NET 343 = spare_buffer_238.q
* NET 358 = spare_buffer_337.q
* NET 360 = m_clock_root_tr_tr_tr_0
* NET 363 = abc_8306_new_n938
* NET 366 = spare_buffer_333.q
* NET 368 = m_clock_root_tr_tr_tl_0
* NET 370 = abc_8306_new_n875
* NET 372 = abc_8306_new_n876
* NET 374 = spare_buffer_321.q
* NET 376 = spare_buffer_320.q
* NET 378 = abc_8306_new_n850
* NET 382 = spare_buffer_317.q
* NET 384 = spare_buffer_316.q
* NET 387 = spare_buffer_257.q
* NET 390 = op_bit5_hfns_2
* NET 392 = spare_buffer_253.q
* NET 396 = spare_buffer_241.q
* NET 399 = abc_8306_new_n335
* NET 401 = spare_buffer_237.q
* NET 403 = m_clock_root_tl_tl_tl_0
* NET 405 = abc_8306_new_n445
* NET 434 = abc_8306_new_n510_hfns_2
* NET 437 = ex_st[1]
* NET 440 = subckt_1575_sff1_x4.sff_m
* NET 443 = subckt_1575_sff1_x4.ckr
* NET 444 = subckt_1575_sff1_x4.nckr
* NET 446 = abc_8306_new_n1303
* NET 455 = abc_8306_new_n916
* NET 461 = abc_8306_new_n873
* NET 462 = abc_8306_new_n877
* NET 464 = abc_8306_new_n775
* NET 468 = abc_8306_new_n783
* NET 469 = abc_8306_new_n781
* NET 470 = abc_8306_new_n777
* NET 478 = subckt_1575_sff1_x4.sff_s
* NET 480 = abc_8306_auto_rtlil_cc_2608_muxgate_8075
* NET 481 = abc_8306_new_n345
* NET 494 = abc_8306_new_n441
* NET 495 = abc_8306_new_n500
* NET 507 = abc_8306_new_n874
* NET 509 = abc_8306_new_n803
* NET 511 = abc_8306_new_n870
* NET 512 = abc_8306_new_n860
* NET 514 = abc_8306_new_n786
* NET 515 = abc_8306_new_n785
* NET 518 = abc_8306_new_n782
* NET 522 = subckt_1612_sff1_x4.sff_s
* NET 526 = subckt_1612_sff1_x4.sff_m
* NET 527 = abc_8306_auto_rtlil_cc_2608_muxgate_8149
* NET 529 = subckt_1612_sff1_x4.ckr
* NET 530 = subckt_1612_sff1_x4.nckr
* NET 533 = abc_8306_new_n436
* NET 536 = abc_8306_new_n438
* NET 554 = abc_8306_new_n937
* NET 558 = abc_8306_new_n940
* NET 563 = abc_8306_new_n827
* NET 564 = abc_8306_new_n867
* NET 566 = abc_8306_new_n866
* NET 568 = abc_8306_new_n859
* NET 571 = abc_8306_new_n861
* NET 576 = abc_8306_new_n778
* NET 579 = op[6]
* NET 580 = subckt_1616_sff1_x4.sff_s
* NET 584 = abc_8306_auto_rtlil_cc_2608_muxgate_8157
* NET 585 = subckt_1616_sff1_x4.sff_m
* NET 587 = subckt_1616_sff1_x4.ckr
* NET 589 = subckt_1616_sff1_x4.nckr
* NET 593 = subckt_1617_sff1_x4.sff_s
* NET 596 = subckt_1617_sff1_x4.sff_m
* NET 598 = m_clock_root_tl_tr_tl_0
* NET 599 = subckt_1617_sff1_x4.ckr
* NET 601 = subckt_1617_sff1_x4.nckr
* NET 602 = ex_st_bit1_hfns_2
* NET 609 = abc_8306_new_n440
* NET 640 = abc_8306_new_n878
* NET 641 = abc_8306_new_n915
* NET 642 = abc_8306_new_n939
* NET 647 = abc_8306_new_n774
* NET 653 = abc_8306_new_n687
* NET 654 = abc_8306_new_n689
* NET 656 = abc_8306_auto_rtlil_cc_2608_muxgate_8155
* NET 662 = subckt_1613_sff1_x4.sff_s
* NET 665 = subckt_1613_sff1_x4.sff_m
* NET 667 = subckt_1613_sff1_x4.ckr
* NET 669 = m_clock_root_tl_tl_tr_0
* NET 670 = subckt_1613_sff1_x4.nckr
* NET 685 = abc_8306_new_n985
* NET 691 = abc_8306_new_n889
* NET 695 = abc_8306_new_n879
* NET 696 = abc_8306_new_n886
* NET 698 = abc_8306_new_n868
* NET 699 = abc_8306_new_n882
* NET 706 = abc_8306_new_n708
* NET 709 = abc_8306_new_n706
* NET 721 = abc_8306_new_n433_hfns_2
* NET 728 = abc_8306_new_n414
* NET 729 = abc_8306_new_n696
* NET 731 = abc_8306_new_n406
* NET 735 = p_reset_hfns_2
* NET 762 = abc_8306_new_n980
* NET 765 = abc_8306_new_n884
* NET 767 = abc_8306_new_n885
* NET 768 = abc_8306_new_n883
* NET 771 = abc_8306_new_n856
* NET 775 = abc_8306_new_n686
* NET 776 = abc_8306_new_n688
* NET 777 = abc_8306_new_n705
* NET 778 = abc_8306_new_n690
* NET 780 = subckt_1614_sff1_x4.sff_s
* NET 784 = subckt_1614_sff1_x4.sff_m
* NET 785 = abc_8306_auto_rtlil_cc_2608_muxgate_8153
* NET 787 = subckt_1614_sff1_x4.ckr
* NET 788 = m_clock_root_tl_tr_tr_0
* NET 789 = subckt_1614_sff1_x4.nckr
* NET 790 = abc_8306_new_n697
* NET 793 = abc_8306_new_n433
* NET 819 = abc_8306_new_n881
* NET 823 = abc_8306_new_n865
* NET 824 = abc_8306_new_n858
* NET 827 = abc_8306_new_n869
* NET 828 = abc_8306_new_n787
* NET 829 = abc_8306_new_n789
* NET 831 = abc_8306_new_n685
* NET 832 = abc_8306_new_n701
* NET 833 = abc_8306_new_n704
* NET 841 = abc_8306_auto_rtlil_cc_2608_muxgate_8151
* NET 844 = abc_8306_new_n348
* NET 847 = abc_8306_new_n501
* NET 875 = abc_8306_new_n449
* NET 890 = abc_8306_new_n1084
* NET 893 = abc_8306_new_n890
* NET 894 = abc_8306_new_n917
* NET 899 = abc_8306_new_n872
* NET 900 = abc_8306_new_n828
* NET 902 = abc_8306_new_n826
* NET 903 = abc_8306_new_n880
* NET 905 = abc_8306_new_n797
* NET 906 = abc_8306_new_n857
* NET 907 = abc_8306_new_n779
* NET 908 = abc_8306_new_n780
* NET 909 = abc_8306_new_n707
* NET 910 = abc_8306_new_n709
* NET 915 = abc_8306_auto_rtlil_cc_2608_muxgate_8159
* NET 918 = abc_8306_new_n357
* NET 936 = abc_8306_new_n991
* NET 937 = abc_8306_new_n989
* NET 939 = abc_8306_new_n975
* NET 942 = abc_8306_new_n981
* NET 949 = abc_8306_new_n795
* NET 951 = abc_8306_new_n669
* NET 953 = abc_8306_new_n710
* NET 960 = abc_8306_new_n703
* NET 963 = tc
* NET 964 = subckt_1666_sff1_x4.sff_s
* NET 968 = abc_8306_auto_rtlil_cc_2608_muxgate_8289
* NET 969 = subckt_1666_sff1_x4.sff_m
* NET 971 = subckt_1666_sff1_x4.ckr
* NET 973 = subckt_1666_sff1_x4.nckr
* NET 975 = abc_8306_new_n698
* NET 978 = abc_8306_new_n430
* NET 979 = abc_8306_new_n432
* NET 1020 = abc_8306_new_n992
* NET 1021 = abc_8306_new_n914
* NET 1022 = abc_8306_new_n988
* NET 1023 = abc_8306_new_n984
* NET 1025 = abc_8306_new_n990
* NET 1029 = abc_8306_new_n887
* NET 1032 = abc_8306_new_n788
* NET 1034 = abc_8306_new_n888
* NET 1037 = abc_8306_new_n683
* NET 1040 = abc_8306_new_n693
* NET 1041 = abc_8306_new_n699
* NET 1044 = abc_8306_new_n609
* NET 1046 = abc_8306_new_n429
* NET 1047 = abc_8306_new_n416
* NET 1049 = abc_8306_new_n344
* NET 1051 = abc_8306_new_n405
* NET 1052 = abc_8306_new_n437
* NET 1068 = abc_8306_new_n974
* NET 1074 = abc_8306_new_n1118
* NET 1075 = abc_8306_new_n1124
* NET 1082 = abc_8306_new_n849
* NET 1085 = abc_8306_new_n672
* NET 1091 = abc_8306_new_n700
* NET 1092 = abc_8306_new_n692
* NET 1106 = abc_8306_new_n431
* NET 1109 = abc_8306_new_n408
* NET 1111 = abc_8306_new_n407
* NET 1112 = abc_8306_new_n415
* NET 1114 = abc_8306_new_n498
* NET 1115 = start
* NET 1144 = abc_8306_new_n1036
* NET 1145 = abc_8306_new_n796
* NET 1146 = abc_8306_new_n1123
* NET 1149 = abc_8306_new_n1121
* NET 1153 = abc_8306_new_n987
* NET 1155 = abc_8306_new_n673
* NET 1159 = abc_8306_new_n1180
* NET 1168 = op[3]
* NET 1180 = spare_buffer_330.q
* NET 1182 = abc_8306_new_n1117
* NET 1185 = spare_buffer_326.q
* NET 1187 = abc_8306_new_n848
* NET 1190 = spare_buffer_314.q
* NET 1196 = spare_buffer_310.q
* NET 1197 = abc_8306_new_n1244
* NET 1201 = spare_buffer_250.q
* NET 1203 = abc_8306_new_n605
* NET 1206 = spare_buffer_246.q
* NET 1210 = spare_buffer_234.q
* NET 1211 = abc_8306_new_n332
* NET 1215 = spare_buffer_230.q
* NET 1216 = abc_8306_new_n1040
* NET 1236 = abc_8306_new_n361
* NET 1253 = spare_buffer_329.q
* NET 1255 = spare_buffer_328.q
* NET 1257 = abc_8306_new_n1041
* NET 1258 = abc_8306_new_n1037
* NET 1261 = spare_buffer_325.q
* NET 1263 = spare_buffer_324.q
* NET 1264 = m_clock_root_tr_tr_0
* NET 1266 = abc_8306_new_n986
* NET 1267 = abc_8306_new_n1242
* NET 1270 = abc_8306_new_n794
* NET 1271 = abc_8306_new_n790
* NET 1273 = spare_buffer_313.q
* NET 1275 = spare_buffer_312.q
* NET 1279 = spare_buffer_309.q
* NET 1282 = spare_buffer_308.q
* NET 1284 = abc_8306_new_n1181
* NET 1287 = abc_8306_new_n900
* NET 1288 = spare_buffer_249.q
* NET 1290 = m_clock_root_tl_tr_br_0
* NET 1292 = abc_8306_new_n435
* NET 1294 = spare_buffer_245.q
* NET 1295 = m_clock_root_tl_tr_0
* NET 1296 = spare_buffer_244.q
* NET 1300 = spare_buffer_233.q
* NET 1302 = spare_buffer_232.q
* NET 1304 = ex_st[4]
* NET 1307 = spare_buffer_229.q
* NET 1309 = spare_buffer_228.q
* NET 1312 = abc_8306_new_n454
* NET 1332 = abc_8306_new_n1093
* NET 1333 = abc_8306_new_n1038
* NET 1334 = abc_8306_new_n1095
* NET 1336 = abc_8306_new_n1101
* NET 1337 = abc_8306_new_n1110
* NET 1339 = abc_8306_new_n1122
* NET 1340 = abc_8306_new_n1120
* NET 1341 = abc_8306_new_n711
* NET 1342 = abc_8306_new_n652
* NET 1355 = abc_8306_new_n750
* NET 1356 = abc_8306_new_n702
* NET 1363 = abc_8306_new_n412
* NET 1365 = abc_8306_new_n359
* NET 1366 = abc_8306_new_n355
* NET 1368 = abc_8306_new_n401
* NET 1369 = abc_8306_new_n598
* NET 1371 = abc_8306_new_n694
* NET 1372 = abc_8306_new_n460
* NET 1373 = abc_8306_new_n695
* NET 1376 = abc_8306_new_n428
* NET 1377 = abc_8306_new_n421
* NET 1382 = abc_8306_new_n497
* NET 1384 = abc_8306_new_n331
* NET 1385 = abc_8306_new_n452
* NET 1412 = p_reset
* NET 1413 = abc_8306_new_n1083
* NET 1419 = abc_8306_new_n1099
* NET 1420 = abc_8306_new_n1098
* NET 1422 = abc_8306_new_n1109
* NET 1426 = abc_8306_new_n1108
* NET 1427 = abc_8306_new_n1058
* NET 1430 = abc_8306_new_n667
* NET 1431 = abc_8306_new_n646
* NET 1435 = abc_8306_new_n645
* NET 1440 = abc_8306_new_n341
* NET 1441 = abc_8306_new_n358
* NET 1444 = abc_8306_new_n458
* NET 1445 = abc_8306_new_n417
* NET 1449 = op[2]
* NET 1464 = abc_8306_new_n1113
* NET 1465 = abc_8306_new_n1114
* NET 1466 = abc_8306_new_n651
* NET 1468 = abc_8306_new_n1111
* NET 1473 = abc_8306_new_n1106
* NET 1474 = abc_8306_new_n1107
* NET 1479 = abc_8306_new_n1102
* NET 1489 = abc_8306_new_n1182
* NET 1496 = abc_8306_new_n721
* NET 1500 = abc_8306_new_n400
* NET 1501 = abc_8306_new_n402
* NET 1508 = abc_8306_new_n484
* NET 1543 = abc_8306_new_n983
* NET 1547 = abc_8306_new_n1126
* NET 1548 = abc_8306_new_n1115
* NET 1550 = abc_8306_new_n1066
* NET 1551 = abc_8306_new_n1100
* NET 1552 = abc_8306_new_n1097
* NET 1556 = abc_8306_new_n1067
* NET 1558 = abc_8306_new_n1064
* NET 1560 = abc_8306_new_n1059
* NET 1565 = abc_8306_new_n1177
* NET 1567 = abc_8306_new_n1176
* NET 1568 = abc_8306_new_n606
* NET 1569 = abc_8306_new_n603
* NET 1570 = abc_8306_new_n600
* NET 1572 = abc_8306_new_n411
* NET 1574 = abc_8306_new_n360
* NET 1575 = abc_8306_new_n342
* NET 1577 = abc_8306_new_n350
* NET 1579 = abc_8306_new_n347
* NET 1581 = abc_8306_new_n424
* NET 1598 = abc_8306_new_n1112
* NET 1605 = abc_8306_new_n1119
* NET 1618 = abc_8306_new_n419
* NET 1619 = abc_8306_new_n404
* NET 1620 = abc_8306_new_n409
* NET 1624 = abc_8306_new_n333
* NET 1627 = abc_8306_new_n496
* NET 1628 = abc_8306_new_n418
* NET 1631 = abc_8306_new_n426
* NET 1632 = abc_8306_new_n499
* NET 1633 = abc_8306_new_n1094
* NET 1634 = abc_8306_new_n1039
* NET 1636 = abc_8306_new_n1096
* NET 1641 = abc_8306_new_n1150
* NET 1652 = abc_8306_new_n607
* NET 1653 = abc_8306_new_n623
* NET 1679 = abc_8306_new_n1032
* NET 1680 = abc_8306_new_n1035
* NET 1681 = abc_8306_new_n1034
* NET 1682 = abc_8306_new_n1105
* NET 1684 = abc_8306_new_n1092
* NET 1686 = abc_8306_new_n1103
* NET 1688 = abc_8306_new_n510_hfns_1
* NET 1694 = abc_8306_new_n1179
* NET 1695 = abc_8306_new_n1178
* NET 1699 = abc_8306_new_n1057
* NET 1700 = abc_8306_new_n653
* NET 1707 = abc_8306_new_n422
* NET 1709 = abc_8306_new_n255
* NET 1723 = abc_8306_new_n1204
* NET 1727 = abc_8306_new_n976
* NET 1728 = abc_8306_new_n982
* NET 1732 = abc_8306_new_n792
* NET 1733 = abc_8306_new_n1169
* NET 1736 = abc_8306_new_n1089
* NET 1740 = abc_8306_new_n1060
* NET 1741 = abc_8306_new_n1065
* NET 1744 = abc_8306_new_n511_hfns_2
* NET 1746 = abc_8306_new_n1794
* NET 1747 = abc_8306_new_n1795
* NET 1749 = abc_8306_new_n1792
* NET 1750 = abc_8306_new_n1793
* NET 1753 = abc_8306_new_n1203
* NET 1759 = abc_8306_new_n553
* NET 1764 = abc_8306_new_n349
* NET 1765 = abc_8306_new_n340
* NET 1767 = abc_8306_new_n648
* NET 1768 = abc_8306_new_n650
* NET 1771 = abc_8306_new_n451
* NET 1775 = abc_8306_new_n336
* NET 1809 = abc_8306_new_n793
* NET 1810 = abc_8306_new_n1116
* NET 1813 = abc_8306_new_n1091
* NET 1819 = abc_8306_new_n1175
* NET 1821 = abc_8306_new_n1174
* NET 1823 = abc_8306_new_n1056
* NET 1825 = abc_8306_new_n746
* NET 1826 = abc_8306_new_n525
* NET 1828 = abc_8306_new_n602
* NET 1830 = abc_8306_new_n610
* NET 1832 = abc_8306_new_n622
* NET 1833 = abc_8306_new_n423
* NET 1834 = abc_8306_new_n550
* NET 1835 = abc_8306_new_n647
* NET 1837 = abc_8306_new_n457
* NET 1838 = abc_8306_new_n448
* NET 1841 = rd
* NET 1851 = abc_8306_new_n684
* NET 1852 = abc_8306_new_n1031
* NET 1855 = abc_8306_new_n1127
* NET 1858 = abc_8306_new_n1043
* NET 1860 = abc_8306_new_n1147
* NET 1866 = abc_8306_new_n668
* NET 1867 = abc_8306_new_n1090
* NET 1869 = abc_8306_new_n1085
* NET 1871 = abc_8306_new_n744
* NET 1872 = abc_8306_new_n751
* NET 1876 = abc_8306_new_n1088
* NET 1880 = abc_8306_new_n551
* NET 1881 = abc_8306_new_n1205
* NET 1883 = abc_8306_new_n1063
* NET 1892 = abc_8306_new_n747
* NET 1893 = abc_8306_new_n636
* NET 1896 = abc_8306_new_n547
* NET 1898 = abc_8306_new_n1202
* NET 1899 = abc_8306_new_n351
* NET 1906 = ex_st[5]
* NET 1908 = abc_8306_new_n346
* NET 1911 = abc_8306_new_n338
* NET 1914 = abc_8306_new_n330
* NET 1915 = abc_8306_new_n329
* NET 1952 = abc_8306_new_n1042
* NET 1954 = abc_8306_new_n1125
* NET 1959 = abc_8306_new_n1082
* NET 1965 = abc_8306_new_n1154
* NET 1967 = abc_8306_new_n1173
* NET 1968 = abc_8306_new_n658
* NET 1970 = abc_8306_new_n627
* NET 1971 = abc_8306_new_n599
* NET 1973 = abc_8306_new_n555
* NET 1974 = abc_8306_new_n560
* NET 1976 = abc_8306_new_n356
* NET 1979 = abc_8306_new_n427
* NET 1981 = rdy_hfns_4
* NET 2002 = abc_8306_new_n1168
* NET 2007 = abc_8306_new_n1149
* NET 2008 = abc_8306_new_n1148
* NET 2009 = abc_8306_new_n1128
* NET 2016 = abc_8306_new_n766
* NET 2018 = abc_8306_new_n752
* NET 2023 = abc_8306_new_n1062
* NET 2027 = abc_8306_new_n1243
* NET 2029 = abc_8306_new_n1245
* NET 2033 = abc_8306_new_n453
* NET 2035 = abc_8306_new_n549
* NET 2037 = abc_8306_new_n554
* NET 2039 = abc_8306_new_n619
* NET 2040 = abc_8306_new_n620
* NET 2041 = abc_8306_new_n621
* NET 2042 = abc_8306_new_n637
* NET 2081 = abc_8306_new_n1167
* NET 2082 = abc_8306_new_n1170
* NET 2085 = abc_8306_new_n995
* NET 2088 = abc_8306_new_n714
* NET 2090 = abc_8306_new_n1157
* NET 2091 = abc_8306_new_n1155
* NET 2093 = abc_8306_new_n1156
* NET 2095 = abc_8306_new_n1080
* NET 2099 = abc_8306_new_n1045
* NET 2101 = abc_8306_new_n1054
* NET 2102 = abc_8306_new_n601
* NET 2103 = abc_8306_new_n248
* NET 2104 = abc_8306_new_n745
* NET 2109 = abc_8306_new_n635
* NET 2111 = op[0]
* NET 2113 = subckt_1610_sff1_x4.sff_s
* NET 2117 = subckt_1610_sff1_x4.sff_m
* NET 2118 = abc_8306_auto_rtlil_cc_2608_muxgate_8145
* NET 2119 = subckt_1610_sff1_x4.ckr
* NET 2121 = subckt_1610_sff1_x4.nckr
* NET 2133 = abc_8306_new_n671
* NET 2134 = abc_8306_new_n824
* NET 2137 = spare_buffer_306.q
* NET 2139 = abc_8306_new_n959
* NET 2140 = abc_8306_new_n996
* NET 2141 = abc_8306_new_n978
* NET 2145 = spare_buffer_302.q
* NET 2149 = abc_8306_new_n921
* NET 2151 = spare_buffer_290.q
* NET 2153 = abc_8306_new_n719
* NET 2154 = abc_8306_new_n718
* NET 2157 = abc_8306_new_n1153
* NET 2159 = abc_8306_new_n1087
* NET 2163 = spare_buffer_286.q
* NET 2164 = abc_8306_new_n715
* NET 2165 = abc_8306_new_n1044
* NET 2168 = abc_8306_new_n626
* NET 2169 = spare_buffer_226.q
* NET 2171 = abc_8306_new_n628
* NET 2174 = abc_8306_new_n459
* NET 2177 = spare_buffer_222.q
* NET 2179 = abc_8306_new_n413
* NET 2182 = abc_8306_new_n630
* NET 2183 = abc_8306_new_n638
* NET 2185 = abc_8306_new_n639
* NET 2187 = spare_buffer_210.q
* NET 2189 = abc_8306_new_n615
* NET 2192 = spare_buffer_206.q
* NET 2213 = spare_buffer_305.q
* NET 2215 = spare_buffer_304.q
* NET 2217 = abc_8306_new_n997
* NET 2220 = abc_8306_new_n722
* NET 2221 = abc_8306_new_n998
* NET 2222 = abc_8306_new_n979
* NET 2224 = spare_buffer_301.q
* NET 2226 = spare_buffer_300.q
* NET 2228 = abc_8306_new_n947
* NET 2229 = abc_8306_new_n894
* NET 2232 = spare_buffer_289.q
* NET 2234 = spare_buffer_288.q
* NET 2237 = spare_buffer_285.q
* NET 2239 = spare_buffer_284.q
* NET 2241 = abc_8306_new_n1055
* NET 2245 = abc_8306_new_n320
* NET 2246 = spare_buffer_225.q
* NET 2252 = spare_buffer_221.q
* NET 2255 = abc_8306_new_n246
* NET 2256 = abc_8306_new_n456
* NET 2257 = abc_8306_new_n545
* NET 2260 = spare_buffer_209.q
* NET 2261 = spare_buffer_208.q
* NET 2263 = abc_8306_new_n569
* NET 2265 = spare_buffer_205.q
* NET 2286 = abc_8306_new_n821
* NET 2287 = abc_8306_new_n822
* NET 2288 = abc_8306_new_n748
* NET 2290 = abc_8306_new_n1027
* NET 2292 = abc_8306_new_n717
* NET 2300 = abc_8306_new_n681
* NET 2304 = abc_8306_new_n1068
* NET 2307 = subckt_1665_sff1_x4.sff_s
* NET 2309 = subckt_1665_sff1_x4.sff_m
* NET 2312 = subckt_1665_sff1_x4.ckr
* NET 2314 = subckt_1665_sff1_x4.nckr
* NET 2315 = abc_8306_new_n530
* NET 2318 = abc_8306_new_n676
* NET 2319 = abc_8306_new_n675
* NET 2322 = abc_8306_new_n425
* NET 2325 = abc_8306_new_n1721
* NET 2328 = abc_8306_new_n633
* NET 2332 = abc_8306_new_n1197
* NET 2333 = abc_8306_new_n1196
* NET 2337 = abc_8306_new_n612
* NET 2338 = abc_8306_new_n557
* NET 2366 = abc_8306_new_n1013
* NET 2371 = abc_8306_new_n855
* NET 2381 = abc_8306_new_n1069
* NET 2383 = abc_8306_new_n1078
* NET 2390 = abc_8306_new_n455
* NET 2392 = abc_8306_new_n353
* NET 2395 = abc_8306_new_n649
* NET 2398 = abc_8306_new_n556
* NET 2412 = abc_8306_new_n818
* NET 2416 = abc_8306_new_n1012
* NET 2418 = abc_8306_new_n960
* NET 2424 = abc_8306_new_n1081
* NET 2425 = abc_8306_new_n898
* NET 2429 = abc_8306_new_n902
* NET 2431 = abc_8306_new_n901
* NET 2433 = abc_8306_new_n682
* NET 2434 = abc_8306_new_n716
* NET 2435 = abc_8306_new_n595
* NET 2442 = abc_8306_new_n321
* NET 2444 = subckt_1611_sff1_x4.sff_s
* NET 2446 = subckt_1611_sff1_x4.sff_m
* NET 2450 = subckt_1611_sff1_x4.ckr
* NET 2451 = subckt_1611_sff1_x4.nckr
* NET 2452 = abc_8306_new_n657
* NET 2454 = abc_8306_new_n487
* NET 2456 = abc_8306_new_n616
* NET 2457 = abc_8306_new_n1742
* NET 2463 = abc_8306_new_n1199
* NET 2465 = abc_8306_new_n1198
* NET 2467 = abc_8306_new_n614
* NET 2502 = abc_8306_new_n749
* NET 2504 = abc_8306_new_n743
* NET 2505 = abc_8306_new_n823
* NET 2507 = abc_8306_new_n1009
* NET 2508 = abc_8306_new_n999
* NET 2510 = abc_8306_new_n772
* NET 2514 = abc_8306_new_n1079
* NET 2517 = abc_8306_new_n315
* NET 2520 = abc_8306_new_n1000
* NET 2521 = abc_8306_new_n948
* NET 2524 = abc_8306_new_n957
* NET 2526 = subckt_1672_sff1r_x4.sff_s
* NET 2529 = subckt_1672_sff1r_x4.sff_m
* NET 2531 = subckt_1672_sff1r_x4.ckr
* NET 2533 = m_clock_root_tl_br_tl_0
* NET 2534 = subckt_1672_sff1r_x4.nckr
* NET 2536 = abc_8306_new_n617
* NET 2537 = abc_8306_new_n489
* NET 2540 = abc_8306_new_n611
* NET 2541 = abc_8306_new_n410
* NET 2542 = abc_8306_new_n420
* NET 2543 = abc_8306_new_n403
* NET 2546 = subckt_1577_sff1_x4.sff_s
* NET 2550 = subckt_1577_sff1_x4.sff_m
* NET 2551 = subckt_1577_sff1_x4.ckr
* NET 2553 = m_clock_root_tl_bl_tl_0
* NET 2554 = subckt_1577_sff1_x4.nckr
* NET 2576 = abc_8306_new_n1030
* NET 2583 = abc_8306_new_n1029
* NET 2587 = abc_8306_new_n1271
* NET 2589 = abc_8306_new_n522
* NET 2590 = abc_8306_new_n316
* NET 2591 = abc_8306_new_n398
* NET 2592 = abc_8306_new_n665
* NET 2596 = ry[7]
* NET 2597 = abc_8306_auto_rtlil_cc_2608_muxgate_8287
* NET 2602 = op[1]
* NET 2603 = abc_8306_auto_rtlil_cc_2608_muxgate_8147
* NET 2608 = abc_8306_new_n1752
* NET 2612 = abc_8306_new_n1753
* NET 2613 = abc_8306_new_n559
* NET 2618 = abc_8306_new_n495
* NET 2620 = abc_8306_new_n488
* NET 2645 = abc_8306_new_n820
* NET 2647 = abc_8306_new_n1134
* NET 2648 = abc_8306_new_n1135
* NET 2652 = abc_8306_new_n1132
* NET 2653 = abc_8306_new_n1131
* NET 2655 = abc_8306_new_n1133
* NET 2657 = abc_8306_new_n724
* NET 2658 = abc_8306_new_n741
* NET 2659 = abc_8306_new_n895
* NET 2661 = abc_8306_new_n739
* NET 2662 = abc_8306_new_n805
* NET 2664 = rx[7]
* NET 2668 = subckt_1657_sff1_x4.sff_s
* NET 2669 = abc_8306_auto_rtlil_cc_2608_muxgate_8271
* NET 2670 = subckt_1657_sff1_x4.sff_m
* NET 2672 = m_clock_root_tl_br_tr_0
* NET 2674 = subckt_1657_sff1_x4.ckr
* NET 2675 = subckt_1657_sff1_x4.nckr
* NET 2676 = abc_8306_new_n529
* NET 2679 = abc_8306_new_n613
* NET 2681 = abc_8306_new_n490
* NET 2684 = abc_8306_new_n558
* NET 2685 = abc_8306_new_n632
* NET 2686 = op_bit5_hfns_1
* NET 2687 = abc_8306_new_n542
* NET 2688 = abc_8306_new_n1785
* NET 2696 = abc_8306_new_n801
* NET 2705 = abc_8306_new_n740
* NET 2707 = abc_8306_new_n893
* NET 2708 = abc_8306_new_n771
* NET 2712 = m_clock_root_tr_0
* NET 2718 = abc_8306_new_n666
* NET 2723 = abc_8306_new_n1053
* NET 2727 = abc_8306_new_n526
* NET 2730 = abc_8306_new_n1722
* NET 2733 = abc_8306_new_n664
* NET 2738 = abc_8306_new_n631
* NET 2739 = abc_8306_new_n662
* NET 2741 = abc_8306_new_n663
* NET 2743 = abc_8306_new_n528
* NET 2746 = m_clock_root_tl_0
* NET 2748 = abc_8306_new_n661
* NET 2751 = abc_8306_new_n1289
* NET 2752 = abc_8306_auto_rtlil_cc_2608_muxgate_8079
* NET 2754 = rdy
* NET 2784 = abc_8306_new_n946
* NET 2785 = abc_8306_new_n817
* NET 2789 = abc_8306_new_n899
* NET 2792 = abc_8306_new_n844
* NET 2794 = abc_8306_new_n742
* NET 2795 = abc_8306_new_n738
* NET 2798 = abc_8306_new_n723
* NET 2800 = abc_8306_new_n643
* NET 2801 = abc_8306_new_n594
* NET 2810 = abc_8306_new_n1077
* NET 2811 = abc_8306_new_n541
* NET 2813 = abc_8306_new_n634
* NET 2814 = abc_8306_new_n544
* NET 2816 = abc_8306_new_n564
* NET 2817 = abc_8306_new_n1256
* NET 2819 = abc_8306_new_n1291
* NET 2820 = abc_8306_new_n1287
* NET 2823 = abc_8306_new_n467
* NET 2825 = abc_8306_new_n1786
* NET 2836 = abc_8306_new_n804
* NET 2837 = abc_8306_new_n815
* NET 2841 = abc_8306_new_n816
* NET 2842 = abc_8306_new_n846
* NET 2844 = abc_8306_new_n897
* NET 2846 = abc_8306_new_n735
* NET 2847 = abc_8306_new_n737
* NET 2853 = abc_8306_new_n644
* NET 2854 = abc_8306_new_n679
* NET 2856 = abc_8306_new_n734
* NET 2860 = abc_8306_new_n1046
* NET 2861 = abc_8306_new_n532
* NET 2862 = abc_8306_new_n593
* NET 2865 = abc_8306_new_n1796
* NET 2866 = abc_8306_auto_rtlil_cc_2608_muxgate_8305
* NET 2869 = abc_8306_new_n1797
* NET 2872 = abc_8306_new_n258
* NET 2875 = abc_8306_new_n1267
* NET 2880 = abc_8306_new_n343
* NET 2881 = abc_8306_new_n247
* NET 2884 = abc_8306_new_n1292
* NET 2887 = abc_8306_new_n1293
* NET 2889 = abc_8306_new_n1301
* NET 2922 = abc_8306_new_n800
* NET 2925 = abc_8306_new_n678
* NET 2926 = abc_8306_new_n656
* NET 2929 = abc_8306_new_n515
* NET 2931 = abc_8306_new_n769
* NET 2932 = abc_8306_new_n1272
* NET 2934 = ry[6]
* NET 2936 = subckt_1664_sff1_x4.sff_s
* NET 2938 = abc_8306_auto_rtlil_cc_2608_muxgate_8285
* NET 2940 = subckt_1664_sff1_x4.sff_m
* NET 2943 = subckt_1664_sff1_x4.ckr
* NET 2944 = subckt_1664_sff1_x4.nckr
* NET 2945 = abc_8306_new_n531
* NET 2946 = abc_8306_new_n524
* NET 2948 = abc_8306_new_n725
* NET 2949 = abc_8306_new_n233
* NET 2951 = abc_8306_new_n1277
* NET 2953 = abc_8306_new_n1791
* NET 2954 = abc_8306_new_n791
* NET 2956 = abc_8306_new_n527
* NET 2958 = abc_8306_new_n674
* NET 2960 = abc_8306_new_n1206
* NET 2963 = subckt_1671_sff1r_x4.sff_s
* NET 2965 = subckt_1671_sff1r_x4.sff_m
* NET 2969 = subckt_1671_sff1r_x4.nckr
* NET 2970 = subckt_1671_sff1r_x4.ckr
* NET 2971 = abc_8306_new_n1787
* NET 2972 = abc_8306_new_n1789
* NET 2973 = abc_8306_auto_rtlil_cc_2608_muxgate_8303
* NET 2986 = abc_8306_new_n1008
* NET 2988 = abc_8306_new_n1193
* NET 2991 = abc_8306_new_n720
* NET 2995 = abc_8306_new_n552
* NET 2999 = abc_8306_new_n1273
* NET 3000 = abc_8306_new_n1086
* NET 3001 = abc_8306_new_n314
* NET 3004 = abc_8306_new_n1061
* NET 3005 = abc_8306_new_n319
* NET 3009 = abc_8306_new_n830
* NET 3012 = abc_8306_new_n234
* NET 3013 = abc_8306_new_n1070
* NET 3023 = abc_8306_new_n486
* NET 3029 = abc_8306_new_n1195
* NET 3030 = abc_8306_new_n1194
* NET 3033 = abc_8306_new_n1200
* NET 3037 = abc_8306_new_n1209
* NET 3066 = abc_8306_new_n944
* NET 3067 = abc_8306_new_n943
* NET 3069 = abc_8306_new_n962
* NET 3070 = abc_8306_new_n963
* NET 3071 = abc_8306_new_n961
* NET 3074 = abc_8306_new_n945
* NET 3077 = abc_8306_new_n839
* NET 3079 = abc_8306_new_n843
* NET 3080 = abc_8306_new_n854
* NET 3081 = abc_8306_new_n511_hfns_1
* NET 3082 = abc_8306_new_n852
* NET 3083 = abc_8306_new_n903
* NET 3084 = abc_8306_new_n896
* NET 3086 = rx[6]
* NET 3088 = subckt_1656_sff1_x4.sff_s
* NET 3091 = subckt_1656_sff1_x4.sff_m
* NET 3092 = abc_8306_auto_rtlil_cc_2608_muxgate_8269
* NET 3095 = subckt_1656_sff1_x4.ckr
* NET 3096 = subckt_1656_sff1_x4.nckr
* NET 3097 = abc_8306_new_n1001
* NET 3100 = subckt_1648_sff1r_x4.sff_s
* NET 3104 = subckt_1648_sff1r_x4.sff_m
* NET 3105 = subckt_1648_sff1r_x4.ckr
* NET 3107 = subckt_1648_sff1r_x4.nckr
* NET 3108 = abc_8306_new_n1799
* NET 3109 = abc_8306_new_n1798
* NET 3116 = abc_8306_new_n1774
* NET 3119 = abc_8306_new_n1208
* NET 3120 = abc_8306_new_n1279
* NET 3128 = abc_8306_new_n814
* NET 3129 = abc_8306_new_n301
* NET 3131 = abc_8306_new_n819
* NET 3132 = spare_buffer_298.q
* NET 3134 = abc_8306_new_n798
* NET 3135 = abc_8306_new_n511_hfns_0
* NET 3137 = abc_8306_new_n840
* NET 3138 = abc_8306_new_n847
* NET 3140 = spare_buffer_294.q
* NET 3142 = abc_8306_new_n922
* NET 3143 = abc_8306_new_n920
* NET 3145 = abc_8306_new_n642
* NET 3147 = spare_buffer_282.q
* NET 3149 = abc_8306_new_n293
* NET 3155 = spare_buffer_278.q
* NET 3156 = abc_8306_new_n813
* NET 3159 = abc_8306_new_n1172
* NET 3160 = abc_8306_new_n1183
* NET 3163 = spare_buffer_218.q
* NET 3167 = abc_8306_new_n510
* NET 3168 = spare_buffer_214.q
* NET 3170 = abc_8306_new_n579
* NET 3176 = spare_buffer_202.q
* NET 3178 = abc_8306_new_n1773
* NET 3179 = abc_8306_new_n1772
* NET 3181 = abc_8306_new_n1777
* NET 3183 = abc_8306_new_n1780
* NET 3184 = abc_8306_new_n1778
* NET 3187 = spare_buffer_198.q
* NET 3204 = spare_buffer_297.q
* NET 3208 = spare_buffer_293.q
* NET 3210 = m_clock_root_tr_br_0
* NET 3212 = abc_8306_new_n625
* NET 3213 = abc_8306_new_n736
* NET 3214 = abc_8306_new_n640
* NET 3216 = abc_8306_new_n1274
* NET 3218 = spare_buffer_281.q
* NET 3220 = spare_buffer_280.q
* NET 3226 = abc_8306_new_n238
* NET 3227 = spare_buffer_277.q
* NET 3232 = abc_8306_new_n733
* NET 3233 = abc_8306_new_n592
* NET 3235 = spare_buffer_217.q
* NET 3238 = abc_8306_new_n949
* NET 3239 = abc_8306_new_n956
* NET 3240 = abc_8306_new_n511
* NET 3244 = spare_buffer_213.q
* NET 3246 = m_clock_root_tl_br_0
* NET 3248 = abc_8306_new_n1286
* NET 3253 = spare_buffer_201.q
* NET 3256 = abc_8306_new_n1213
* NET 3259 = abc_8306_new_n1788
* NET 3261 = spare_buffer_197.q
* NET 3263 = m_clock_root_tl_bl_bl_0
* NET 3264 = m_clock_root_tl_bl_0
* NET 3266 = abc_8306_new_n472
* NET 3287 = subckt_1660_sff1_x4.sff_s
* NET 3290 = subckt_1660_sff1_x4.sff_m
* NET 3294 = subckt_1660_sff1_x4.ckr
* NET 3295 = subckt_1660_sff1_x4.nckr
* NET 3300 = abc_8306_new_n929
* NET 3303 = abc_8306_new_n1276
* NET 3304 = abc_8306_new_n1275
* NET 3311 = subckt_1647_sff1r_x4.sff_s
* NET 3314 = subckt_1647_sff1r_x4.sff_m
* NET 3315 = abc_8306_auto_rtlil_cc_2608_muxgate_8243
* NET 3318 = subckt_1647_sff1r_x4.nckr
* NET 3319 = subckt_1647_sff1r_x4.ckr
* NET 3321 = abc_8306_new_n806
* NET 3322 = abc_8306_new_n548
* NET 3324 = abc_8306_auto_rtlil_cc_2608_muxgate_8249
* NET 3326 = abc_8306_new_n1159
* NET 3334 = subckt_1569_sff1r_x4.sff_s
* NET 3337 = subckt_1569_sff1r_x4.sff_m
* NET 3338 = abc_8306_auto_rtlil_cc_2608_muxgate_8063
* NET 3341 = subckt_1569_sff1r_x4.nckr
* NET 3342 = subckt_1569_sff1r_x4.ckr
* NET 3343 = abc_8306_new_n1249
* NET 3346 = abc_8306_new_n1268
* NET 3347 = abc_8306_new_n1257
* NET 3348 = abc_8306_new_n1255
* NET 3351 = abc_8306_new_n1776
* NET 3352 = op_bit6_hfns_1
* NET 3356 = abc_8306_new_n1779
* NET 3387 = abc_8306_new_n1185
* NET 3389 = abc_8306_new_n1186
* NET 3394 = subckt_1652_sff1_x4.sff_s
* NET 3397 = subckt_1652_sff1_x4.sff_m
* NET 3400 = m_clock_root_tr_br_br_0
* NET 3401 = subckt_1652_sff1_x4.ckr
* NET 3402 = subckt_1652_sff1_x4.nckr
* NET 3403 = abc_8306_new_n842
* NET 3406 = abc_8306_new_n924
* NET 3407 = abc_8306_new_n925
* NET 3409 = abc_8306_new_n919
* NET 3410 = abc_8306_new_n1138
* NET 3411 = abc_8306_new_n1136
* NET 3412 = abc_8306_new_n1130
* NET 3418 = abc_8306_new_n521
* NET 3420 = abc_8306_new_n654
* NET 3422 = subckt_335_nmx2_x1.q
* NET 3425 = abc_8306_new_n399
* NET 3427 = abc_8306_new_n259
* NET 3428 = abc_8306_new_n354
* NET 3431 = abc_8306_new_n482
* NET 3432 = abc_8306_new_n481
* NET 3455 = subckt_1640_sff1_x4.sff_m
* NET 3456 = abc_8306_new_n618
* NET 3462 = subckt_1669_sff1r_x4.sff_m
* NET 3463 = abc_8306_auto_rtlil_cc_2608_muxgate_8299
* NET 3466 = m_clock_root_tl_bl_br_0
* NET 3467 = subckt_1669_sff1r_x4.nckr
* NET 3468 = subckt_1669_sff1r_x4.ckr
* NET 3469 = abc_8306_new_n994
* NET 3470 = abc_8306_new_n993
* NET 3472 = abc_8306_new_n1014
* NET 3475 = ry[2]
* NET 3476 = abc_8306_auto_rtlil_cc_2608_muxgate_8277
* NET 3481 = abc_8306_new_n297
* NET 3482 = abc_8306_new_n845
* NET 3483 = abc_8306_new_n829
* NET 3484 = abc_8306_new_n841
* NET 3487 = abc_8306_new_n927
* NET 3495 = abc_8306_new_n906
* NET 3499 = abc_8306_new_n235
* NET 3500 = abc_8306_new_n239
* NET 3501 = abc_8306_new_n546
* NET 3502 = abc_8306_new_n726
* NET 3504 = subckt_1640_sff1_x4.sff_s
* NET 3507 = subckt_1640_sff1_x4.ckr
* NET 3508 = subckt_1640_sff1_x4.nckr
* NET 3511 = subckt_1669_sff1r_x4.sff_s
* NET 3513 = abc_8306_new_n1212
* NET 3515 = abc_8306_new_n1775
* NET 3516 = abc_8306_new_n1269
* NET 3545 = abc_8306_new_n670
* NET 3546 = abc_8306_new_n510_hfns_0
* NET 3548 = abc_8306_new_n1026
* NET 3549 = abc_8306_new_n1011
* NET 3550 = ry[1]
* NET 3552 = subckt_1659_sff1_x4.sff_s
* NET 3554 = abc_8306_auto_rtlil_cc_2608_muxgate_8275
* NET 3556 = subckt_1659_sff1_x4.sff_m
* NET 3558 = m_clock_root_tr_br_bl_0
* NET 3560 = subckt_1659_sff1_x4.ckr
* NET 3561 = subckt_1659_sff1_x4.nckr
* NET 3562 = abc_8306_new_n926
* NET 3563 = abc_8306_new_n923
* NET 3565 = subckt_1644_sff1r_x4.sff_s
* NET 3568 = abc_8306_auto_rtlil_cc_2608_muxgate_8225
* NET 3570 = subckt_1644_sff1r_x4.sff_m
* NET 3571 = m_clock_root_tr_bl_bl_0
* NET 3572 = subckt_1644_sff1r_x4.ckr
* NET 3574 = subckt_1644_sff1r_x4.nckr
* NET 3576 = subckt_1649_sff1r_x4.sff_s
* NET 3579 = subckt_1649_sff1r_x4.sff_m
* NET 3581 = m_clock_root_tl_br_br_0
* NET 3582 = abc_8306_auto_rtlil_cc_2608_muxgate_8255
* NET 3583 = subckt_1649_sff1r_x4.ckr
* NET 3585 = subckt_1649_sff1r_x4.nckr
* NET 3586 = subckt_1641_sff1_x4.sff_s
* NET 3590 = subckt_1641_sff1_x4.sff_m
* NET 3592 = abc_8306_auto_rtlil_cc_2608_muxgate_8207
* NET 3594 = subckt_1641_sff1_x4.ckr
* NET 3595 = m_clock_root_tl_br_bl_0
* NET 3596 = subckt_1641_sff1_x4.nckr
* NET 3601 = abc_8306_new_n1767
* NET 3625 = abc_8306_new_n1028
* NET 3632 = abc_8306_new_n942
* NET 3633 = abc_8306_new_n964
* NET 3636 = abc_8306_new_n904
* NET 3637 = abc_8306_new_n892
* NET 3644 = abc_8306_new_n237
* NET 3645 = abc_8306_new_n240
* NET 3646 = abc_8306_new_n236
* NET 3648 = abc_8306_auto_rtlil_cc_2608_muxgate_8205
* NET 3649 = abc_8306_new_n1160
* NET 3655 = abc_8306_new_n1246
* NET 3659 = abc_8306_new_n1254
* NET 3660 = abc_8306_new_n1253
* NET 3663 = abc_8306_new_n1201
* NET 3665 = abc_8306_new_n257
* NET 3666 = abc_8306_new_n1770
* NET 3667 = abc_8306_new_n1210
* NET 3670 = abc_8306_new_n475
* NET 3695 = abc_8306_auto_rtlil_cc_2608_muxgate_8261
* NET 3696 = rx[2]
* NET 3701 = abc_8306_new_n853
* NET 3705 = abc_8306_new_n296
* NET 3710 = abc_8306_new_n289
* NET 3713 = abc_8306_new_n755
* NET 3717 = m_clock
* NET 3719 = abc_8306_new_n831
* NET 3720 = abc_8306_new_n838
* NET 3722 = abc_8306_new_n812
* NET 3724 = abc_8306_new_n273
* NET 3727 = ra[6]
* NET 3729 = abc_8306_new_n1732
* NET 3732 = abc_8306_new_n562
* NET 3733 = abc_8306_new_n563
* NET 3734 = abc_8306_new_n568
* NET 3736 = abc_8306_new_n1782
* NET 3737 = abc_8306_new_n1783
* NET 3738 = abc_8306_new_n1211
* NET 3739 = abc_8306_new_n260
* NET 3742 = abc_8306_new_n251
* NET 3743 = abc_8306_new_n1768
* NET 3744 = abc_8306_new_n1337
* NET 3769 = abc_8306_new_n1010
* NET 3770 = abc_8306_new_n311
* NET 3771 = abc_8306_new_n310
* NET 3774 = rx[1]
* NET 3776 = subckt_1651_sff1_x4.sff_s
* NET 3779 = abc_8306_auto_rtlil_cc_2608_muxgate_8259
* NET 3780 = subckt_1651_sff1_x4.sff_m
* NET 3782 = subckt_1651_sff1_x4.ckr
* NET 3784 = subckt_1651_sff1_x4.nckr
* NET 3791 = subckt_1643_sff1r_x4.sff_s
* NET 3795 = subckt_1643_sff1r_x4.sff_m
* NET 3797 = abc_8306_auto_rtlil_cc_2608_muxgate_8219
* NET 3799 = subckt_1643_sff1r_x4.ckr
* NET 3800 = subckt_1643_sff1r_x4.nckr
* NET 3804 = abc_8306_new_n930
* NET 3810 = abc_8306_new_n1076
* NET 3811 = abc_8306_new_n284
* NET 3814 = fd
* NET 3817 = abc_8306_new_n566
* NET 3819 = fv
* NET 3820 = op[7]
* NET 3827 = subckt_1670_sff1r_x4.sff_s
* NET 3830 = abc_8306_auto_rtlil_cc_2608_muxgate_8301
* NET 3831 = subckt_1670_sff1r_x4.sff_m
* NET 3834 = subckt_1670_sff1r_x4.ckr
* NET 3835 = subckt_1670_sff1r_x4.nckr
* NET 3836 = abc_8306_new_n1769
* NET 3837 = abc_8306_new_n565
* NET 3840 = abc_8306_new_n538
* NET 3868 = rx[3]
* NET 3870 = abc_8306_new_n967
* NET 3876 = abc_8306_auto_rtlil_cc_2608_muxgate_8263
* NET 3878 = abc_8306_new_n799
* NET 3879 = ry[0]
* NET 3881 = subckt_1658_sff1_x4.sff_s
* NET 3884 = abc_8306_auto_rtlil_cc_2608_muxgate_8273
* NET 3885 = subckt_1658_sff1_x4.sff_m
* NET 3888 = subckt_1658_sff1_x4.nckr
* NET 3889 = subckt_1658_sff1_x4.ckr
* NET 3890 = ra[3]
* NET 3893 = subckt_1637_sff1_x4.sff_s
* NET 3895 = abc_8306_auto_rtlil_cc_2608_muxgate_8199
* NET 3896 = subckt_1637_sff1_x4.sff_m
* NET 3899 = subckt_1637_sff1_x4.ckr
* NET 3900 = subckt_1637_sff1_x4.nckr
* NET 3902 = subckt_1646_sff1r_x4.sff_s
* NET 3905 = abc_8306_auto_rtlil_cc_2608_muxgate_8237
* NET 3907 = subckt_1646_sff1r_x4.sff_m
* NET 3909 = subckt_1646_sff1r_x4.nckr
* NET 3910 = subckt_1646_sff1r_x4.ckr
* NET 3911 = abc_8306_new_n1052
* NET 3913 = abc_8306_new_n287
* NET 3917 = abc_8306_new_n1247
* NET 3920 = abc_8306_new_n573
* NET 3922 = abc_8306_new_n1207
* NET 3925 = abc_8306_new_n471
* NET 3927 = abc_8306_new_n537
* NET 3951 = subckt_1642_sff1r_x4.sff_m
* NET 3953 = abc_8306_auto_rtlil_cc_2608_muxgate_8213
* NET 3955 = subckt_1642_sff1r_x4.ckr
* NET 3956 = subckt_1642_sff1r_x4.nckr
* NET 3957 = abc_8306_new_n753
* NET 3958 = abc_8306_new_n712
* NET 3961 = subckt_1635_sff1_x4.sff_m
* NET 3966 = abc_8306_new_n567
* NET 3967 = abc_8306_new_n571
* NET 3978 = abc_8306_new_n309
* NET 3979 = abc_8306_new_n977
* NET 3982 = subckt_1642_sff1r_x4.sff_s
* NET 3984 = subckt_1635_sff1_x4.sff_s
* NET 3986 = subckt_1635_sff1_x4.ckr
* NET 3988 = subckt_1635_sff1_x4.nckr
* NET 3989 = abc_8306_new_n732
* NET 3992 = abc_8306_new_n267
* NET 3993 = fz
* NET 3997 = ra[7]
* NET 4000 = abc_8306_new_n249
* NET 4006 = abc_8306_new_n1252
* NET 4037 = subckt_1620_sff1_x4.sff_s
* NET 4040 = abc_8306_auto_rtlil_cc_2608_muxgate_8165
* NET 4042 = subckt_1620_sff1_x4.sff_m
* NET 4044 = subckt_1620_sff1_x4.nckr
* NET 4045 = subckt_1620_sff1_x4.ckr
* NET 4047 = subckt_1645_sff1r_x4.sff_s
* NET 4048 = subckt_1645_sff1r_x4.sff_m
* NET 4053 = subckt_1645_sff1r_x4.nckr
* NET 4054 = subckt_1645_sff1r_x4.ckr
* NET 4057 = subckt_1636_sff1_x4.sff_s
* NET 4059 = abc_8306_auto_rtlil_cc_2608_muxgate_8197
* NET 4060 = subckt_1636_sff1_x4.sff_m
* NET 4063 = subckt_1636_sff1_x4.ckr
* NET 4064 = subckt_1636_sff1_x4.nckr
* NET 4066 = abc_8306_new_n591
* NET 4067 = abc_8306_new_n265
* NET 4069 = ra[2]
* NET 4070 = abc_8306_new_n955
* NET 4074 = abc_8306_new_n1248
* NET 4075 = abc_8306_new_n1346
* NET 4077 = abc_8306_new_n574
* NET 4079 = abc_8306_new_n570
* NET 4081 = abc_8306_new_n433_hfns_1
* NET 4084 = abc_8306_new_n1251
* NET 4103 = abc_8306_auto_rtlil_cc_2608_muxgate_8265
* NET 4104 = rx[4]
* NET 4106 = abc_8306_new_n1743
* NET 4112 = abc_8306_new_n304
* NET 4113 = rx[0]
* NET 4115 = subckt_1650_sff1_x4.sff_s
* NET 4118 = subckt_1650_sff1_x4.sff_m
* NET 4119 = abc_8306_auto_rtlil_cc_2608_muxgate_8257
* NET 4122 = subckt_1650_sff1_x4.nckr
* NET 4123 = subckt_1650_sff1_x4.ckr
* NET 4124 = subckt_1634_sff1_x4.sff_s
* NET 4128 = subckt_1634_sff1_x4.sff_m
* NET 4131 = subckt_1634_sff1_x4.nckr
* NET 4132 = subckt_1634_sff1_x4.ckr
* NET 4134 = subckt_1639_sff1_x4.sff_s
* NET 4136 = subckt_1639_sff1_x4.sff_m
* NET 4140 = subckt_1639_sff1_x4.ckr
* NET 4141 = subckt_1639_sff1_x4.nckr
* NET 4142 = abc_8306_new_n837
* NET 4143 = abc_8306_new_n270
* NET 4148 = fc
* NET 4149 = abc_8306_new_n761
* NET 4156 = fn
* NET 4157 = abc_8306_new_n572
* NET 4158 = op_bit5_hfns_0
* NET 4161 = op[4]
* NET 4166 = subckt_1668_sff1r_x4.sff_s
* NET 4170 = subckt_1668_sff1r_x4.sff_m
* NET 4172 = abc_8306_auto_rtlil_cc_2608_muxgate_8297
* NET 4173 = subckt_1668_sff1r_x4.ckr
* NET 4175 = subckt_1668_sff1r_x4.nckr
* NET 4193 = spare_buffer_178.q
* NET 4195 = abc_8306_new_n1609
* NET 4197 = abc_8306_new_n300
* NET 4198 = spare_buffer_174.q
* NET 4204 = spare_buffer_162.q
* NET 4206 = abc_8306_auto_rtlil_cc_2608_muxgate_8193
* NET 4207 = ra[0]
* NET 4211 = abc_8306_new_n756
* NET 4213 = spare_buffer_158.q
* NET 4215 = ra[1]
* NET 4216 = abc_8306_auto_rtlil_cc_2608_muxgate_8195
* NET 4217 = abc_8306_new_n907
* NET 4222 = spare_buffer_98.q
* NET 4224 = abc_8306_new_n514
* NET 4226 = spare_buffer_94.q
* NET 4228 = abc_8306_new_n759
* NET 4231 = abc_8306_new_n1654
* NET 4232 = spare_buffer_82.q
* NET 4236 = spare_buffer_78.q
* NET 4245 = spare_buffer_177.q
* NET 4247 = spare_buffer_176.q
* NET 4249 = abc_8306_new_n1622
* NET 4251 = spare_buffer_173.q
* NET 4254 = abc_8306_new_n770
* NET 4255 = abc_8306_new_n292
* NET 4258 = spare_buffer_161.q
* NET 4261 = abc_8306_auto_rtlil_cc_2608_muxgate_8231
* NET 4264 = abc_8306_new_n1733
* NET 4265 = abc_8306_new_n966
* NET 4268 = spare_buffer_157.q
* NET 4275 = spare_buffer_97.q
* NET 4277 = m_clock_root_bl_tr_tr_0
* NET 4282 = abc_8306_new_n278
* NET 4283 = spare_buffer_93.q
* NET 4292 = spare_buffer_81.q
* NET 4294 = spare_buffer_80.q
* NET 4296 = abc_8306_new_n1290
* NET 4297 = abc_8306_new_n1653
* NET 4303 = spare_buffer_77.q
* NET 4305 = m_clock_root_bl_tl_tl_0
* NET 4339 = subckt_1622_sff1_x4.sff_s
* NET 4342 = subckt_1622_sff1_x4.sff_m
* NET 4345 = subckt_1622_sff1_x4.ckr
* NET 4346 = subckt_1622_sff1_x4.nckr
* NET 4347 = subckt_1625_sff1_x4.sff_s
* NET 4352 = subckt_1625_sff1_x4.sff_m
* NET 4354 = subckt_1625_sff1_x4.ckr
* NET 4355 = subckt_1625_sff1_x4.nckr
* NET 4359 = abc_8306_new_n1007
* NET 4360 = abc_8306_new_n561
* NET 4361 = abc_8306_new_n281
* NET 4364 = abc_8306_new_n1655
* NET 4367 = abc_8306_new_n517
* NET 4368 = abc_8306_new_n518
* NET 4370 = abc_8306_new_n1260
* NET 4372 = abc_8306_new_n1266
* NET 4376 = ex
* NET 4377 = abc_8306_new_n373
* NET 4378 = abc_8306_new_n232
* NET 4395 = subckt_1602_sff1_x4.sff_m
* NET 4401 = abc_8306_new_n1581
* NET 4405 = subckt_1602_sff1_x4.sff_s
* NET 4408 = subckt_1602_sff1_x4.nckr
* NET 4409 = subckt_1602_sff1_x4.ckr
* NET 4410 = abc_8306_new_n680
* NET 4411 = abc_8306_new_n655
* NET 4412 = abc_8306_new_n288
* NET 4413 = abc_8306_new_n677
* NET 4416 = abc_8306_auto_rtlil_cc_2608_muxgate_8175
* NET 4424 = abc_8306_auto_ff_cc_704_flip_bits_8244
* NET 4425 = abc_8306_new_n1563
* NET 4427 = abc_8306_new_n1458
* NET 4431 = abc_8306_auto_ff_cc_704_flip_bits_8208
* NET 4437 = abc_8306_new_n397
* NET 4441 = abc_8306_new_n379
* NET 4442 = abc_8306_new_n372
* NET 4446 = abc_8306_new_n334
* NET 4447 = abc_8306_new_n374
* NET 4448 = abc_8306_new_n378
* NET 4474 = subckt_1623_sff1_x4.sff_s
* NET 4475 = abc_8306_auto_rtlil_cc_2608_muxgate_8171
* NET 4477 = subckt_1623_sff1_x4.sff_m
* NET 4480 = subckt_1623_sff1_x4.ckr
* NET 4481 = subckt_1623_sff1_x4.nckr
* NET 4484 = subckt_1618_sff1_x4.sff_s
* NET 4486 = subckt_1618_sff1_x4.sff_m
* NET 4488 = m_clock_root_br_tl_tr_0
* NET 4490 = subckt_1618_sff1_x4.ckr
* NET 4491 = subckt_1618_sff1_x4.nckr
* NET 4493 = subckt_1638_sff1_x4.sff_s
* NET 4497 = subckt_1638_sff1_x4.sff_m
* NET 4498 = abc_8306_auto_rtlil_cc_2608_muxgate_8201
* NET 4500 = subckt_1638_sff1_x4.ckr
* NET 4501 = subckt_1638_sff1_x4.nckr
* NET 4502 = abc_8306_auto_ff_cc_704_flip_bits_8238
* NET 4504 = abc_8306_auto_ff_cc_704_flip_bits_8250
* NET 4511 = abc_8306_new_n596
* NET 4514 = abc_8306_new_n1265
* NET 4517 = abc_8306_new_n450
* NET 4518 = abc_8306_new_n442
* NET 4524 = abc_8306_new_n494
* NET 4541 = subckt_1603_sff1_x4.sff_s
* NET 4545 = subckt_1603_sff1_x4.sff_m
* NET 4548 = subckt_1603_sff1_x4.nckr
* NET 4549 = subckt_1603_sff1_x4.ckr
* NET 4555 = subckt_1624_sff1_x4.sff_s
* NET 4557 = subckt_1624_sff1_x4.sff_m
* NET 4561 = m_clock_root_br_tl_tl_0
* NET 4562 = subckt_1624_sff1_x4.ckr
* NET 4563 = subckt_1624_sff1_x4.nckr
* NET 4566 = abc_8306_new_n520
* NET 4568 = abc_8306_new_n629
* NET 4569 = abc_8306_new_n604
* NET 4572 = abc_8306_auto_rtlil_cc_2608_muxgate_8203
* NET 4574 = abc_8306_new_n1139
* NET 4577 = abc_8306_new_n1723
* NET 4579 = abc_8306_new_n1461
* NET 4581 = abc_8306_new_n1463
* NET 4582 = abc_8306_new_n1460
* NET 4583 = abc_8306_new_n691
* NET 4585 = abc_8306_new_n1462
* NET 4588 = abc_8306_new_n608
* NET 4589 = abc_8306_new_n580
* NET 4593 = abc_8306_new_n253
* NET 4594 = abc_8306_new_n381
* NET 4597 = abc_8306_new_n339
* NET 4600 = abc_8306_new_n433_hfns_0
* NET 4602 = abc_8306_new_n447
* NET 4603 = abc_8306_new_n446
* NET 4604 = abc_8306_new_n493
* NET 4629 = abc_8306_new_n1620
* NET 4630 = subckt_1621_sff1_x4.sff_s
* NET 4633 = subckt_1621_sff1_x4.sff_m
* NET 4635 = abc_8306_auto_rtlil_cc_2608_muxgate_8167
* NET 4638 = m_clock_root_br_tr_tl_0
* NET 4639 = subckt_1621_sff1_x4.ckr
* NET 4640 = subckt_1621_sff1_x4.nckr
* NET 4641 = abc_8306_auto_rtlil_cc_2608_muxgate_8131
* NET 4642 = adrs[8]
* NET 4644 = abc_8306_auto_rtlil_cc_2608_muxgate_8173
* NET 4649 = abc_8306_new_n1550
* NET 4651 = abc_8306_new_n1576
* NET 4654 = subckt_1598_sff1_x4.sff_s
* NET 4658 = subckt_1598_sff1_x4.sff_m
* NET 4660 = m_clock_root_bl_tr_tl_0
* NET 4661 = subckt_1598_sff1_x4.ckr
* NET 4662 = subckt_1598_sff1_x4.nckr
* NET 4667 = abc_8306_new_n660
* NET 4669 = abc_8306_new_n540
* NET 4673 = abc_8306_new_n1336
* NET 4674 = abc_8306_new_n543
* NET 4676 = abc_8306_new_n492
* NET 4679 = abc_8306_new_n470
* NET 4694 = abc_8306_new_n958
* NET 4695 = abc_8306_new_n624
* NET 4696 = abc_8306_new_n306
* NET 4697 = abc_8306_new_n641
* NET 4698 = abc_8306_new_n305
* NET 4701 = abc_8306_new_n1623
* NET 4702 = abc_8306_new_n1627
* NET 4705 = abc_8306_auto_rtlil_cc_2608_muxgate_8169
* NET 4710 = abc_8306_auto_rtlil_cc_2608_muxgate_8161
* NET 4715 = abc_8306_new_n1590
* NET 4716 = abc_8306_auto_ff_cc_704_flip_bits_8226
* NET 4718 = abc_8306_auto_ff_cc_704_flip_bits_8232
* NET 4720 = abc_8306_new_n1555
* NET 4722 = abc_8306_new_n1537
* NET 4724 = abc_8306_new_n513
* NET 4726 = abc_8306_new_n523
* NET 4728 = abc_8306_new_n439
* NET 4732 = abc_8306_new_n539
* NET 4752 = abc_8306_new_n1619
* NET 4754 = abc_8306_new_n1613
* NET 4755 = abc_8306_new_n1610
* NET 4758 = abc_8306_new_n1614
* NET 4760 = abc_8306_new_n1600
* NET 4762 = abc_8306_new_n1595
* NET 4764 = abc_8306_new_n1583
* NET 4765 = abc_8306_auto_rtlil_cc_2608_muxgate_8129
* NET 4769 = abc_8306_new_n1525
* NET 4771 = abc_8306_new_n1564
* NET 4773 = abc_8306_new_n597
* NET 4774 = abc_8306_new_n1589
* NET 4777 = abc_8306_new_n1466
* NET 4779 = abc_8306_auto_rtlil_cc_2608_muxgate_8121
* NET 4780 = abc_8306_new_n1283
* NET 4781 = abc_8306_new_n519
* NET 4782 = ra[4]
* NET 4783 = abc_8306_new_n505
* NET 4789 = abc_8306_new_n462
* NET 4790 = abc_8306_new_n491
* NET 4809 = abc_8306_new_n1629
* NET 4813 = subckt_1600_sff1_x4.sff_m
* NET 4815 = abc_8306_new_n507
* NET 4819 = abc_8306_new_n1465
* NET 4820 = abc_8306_new_n1459
* NET 4821 = abc_8306_new_n1464
* NET 4822 = abc_8306_new_n1284
* NET 4823 = abc_8306_new_n1285
* NET 4824 = abc_8306_new_n1324
* NET 4825 = abc_8306_new_n1345
* NET 4827 = abc_8306_new_n1264
* NET 4828 = abc_8306_new_n533
* NET 4829 = abc_8306_new_n534
* NET 4833 = abc_8306_new_n1616
* NET 4834 = data[4]
* NET 4837 = abc_8306_new_n1618
* NET 4838 = abc_8306_new_n313
* NET 4841 = abc_8306_new_n295
* NET 4846 = abc_8306_new_n1593
* NET 4847 = abc_8306_new_n1592
* NET 4848 = abc_8306_new_n1586
* NET 4852 = abc_8306_new_n318
* NET 4855 = subckt_1600_sff1_x4.sff_s
* NET 4857 = abc_8306_auto_rtlil_cc_2608_muxgate_8125
* NET 4859 = subckt_1600_sff1_x4.ckr
* NET 4860 = subckt_1600_sff1_x4.nckr
* NET 4861 = abc_8306_auto_ff_cc_704_flip_bits_8214
* NET 4862 = abc_8306_new_n1495
* NET 4869 = abc_8306_new_n480
* NET 4899 = subckt_1604_sff1_x4.sff_s
* NET 4903 = subckt_1604_sff1_x4.sff_m
* NET 4904 = subckt_1604_sff1_x4.ckr
* NET 4906 = subckt_1604_sff1_x4.nckr
* NET 4908 = abc_8306_new_n303
* NET 4912 = abc_8306_new_n1656
* NET 4916 = abc_8306_new_n291
* NET 4920 = abc_8306_new_n1551
* NET 4921 = abc_8306_new_n1549
* NET 4923 = abc_8306_new_n1562
* NET 4926 = abc_8306_new_n1536
* NET 4927 = abc_8306_new_n1538
* NET 4929 = abc_8306_new_n1479
* NET 4933 = ra[5]
* NET 4934 = op_bit6_hfns_0
* NET 4937 = abc_8306_auto_ff_cc_704_flip_bits_8292
* NET 4938 = irq
* NET 4959 = adrs[11]
* NET 4961 = subckt_1605_sff1_x4.sff_s
* NET 4963 = subckt_1605_sff1_x4.sff_m
* NET 4966 = abc_8306_auto_rtlil_cc_2608_muxgate_8135
* NET 4967 = subckt_1605_sff1_x4.ckr
* NET 4969 = subckt_1605_sff1_x4.nckr
* NET 4971 = abc_8306_new_n299
* NET 4973 = abc_8306_new_n1599
* NET 4975 = adrs[9]
* NET 4978 = abc_8306_new_n1596
* NET 4979 = data[6]
* NET 4982 = abc_8306_new_n1634
* NET 4984 = abc_8306_new_n1152
* NET 4985 = abc_8306_new_n516
* NET 4986 = abc_8306_new_n1158
* NET 4987 = abc_8306_new_n1151
* NET 4991 = abc_8306_auto_ff_cc_704_flip_bits_8220
* NET 4995 = abc_8306_new_n1281
* NET 4996 = abc_8306_new_n1280
* NET 4998 = abc_8306_new_n1161
* NET 5000 = abc_8306_new_n250
* NET 5001 = ex_st_bit1_hfns_1
* NET 5006 = subckt_1585_sff1r_x4.sff_s
* NET 5010 = subckt_1585_sff1r_x4.sff_m
* NET 5012 = abc_8306_auto_rtlil_cc_2608_muxgate_8095
* NET 5013 = subckt_1585_sff1r_x4.ckr
* NET 5015 = subckt_1585_sff1r_x4.nckr
* NET 5016 = abc_8306_new_n483
* NET 5043 = data[0]
* NET 5045 = adrs[12]
* NET 5046 = subckt_1606_sff1_x4.sff_s
* NET 5050 = subckt_1606_sff1_x4.sff_m
* NET 5051 = abc_8306_auto_rtlil_cc_2608_muxgate_8137
* NET 5053 = subckt_1606_sff1_x4.ckr
* NET 5054 = subckt_1606_sff1_x4.nckr
* NET 5055 = data[1]
* NET 5056 = abc_8306_new_n1598
* NET 5060 = subckt_1619_sff1_x4.sff_s
* NET 5064 = subckt_1619_sff1_x4.sff_m
* NET 5065 = abc_8306_auto_rtlil_cc_2608_muxgate_8163
* NET 5067 = subckt_1619_sff1_x4.ckr
* NET 5068 = subckt_1619_sff1_x4.nckr
* NET 5069 = abc_8306_new_n1582
* NET 5071 = abc_8306_new_n1588
* NET 5072 = abc_8306_new_n1587
* NET 5074 = abc_8306_new_n1526
* NET 5075 = abc_8306_new_n1523
* NET 5078 = abc_8306_new_n1566
* NET 5079 = abc_8306_new_n1565
* NET 5082 = abc_8306_new_n1478
* NET 5083 = abc_8306_new_n1480
* NET 5085 = abc_8306_new_n584
* NET 5087 = abc_8306_new_n1473
* NET 5092 = abc_8306_new_n1326
* NET 5093 = abc_8306_new_n659
* NET 5097 = abc_8306_new_n1263
* NET 5099 = subckt_1570_sff1r_x4.sff_s
* NET 5100 = p_reset_hfns_1
* NET 5103 = subckt_1570_sff1r_x4.sff_m
* NET 5106 = subckt_1570_sff1r_x4.ckr
* NET 5107 = subckt_1570_sff1r_x4.nckr
* NET 5124 = abc_8306_auto_rtlil_cc_2608_muxgate_8281
* NET 5125 = ry[4]
* NET 5127 = abc_8306_new_n1016
* NET 5128 = abc_8306_new_n1754
* NET 5134 = abc_8306_new_n308
* NET 5137 = data[5]
* NET 5138 = data[7]
* NET 5141 = subckt_1601_sff1_x4.sff_s
* NET 5144 = subckt_1601_sff1_x4.sff_m
* NET 5148 = subckt_1601_sff1_x4.ckr
* NET 5149 = subckt_1601_sff1_x4.nckr
* NET 5153 = abc_8306_new_n1511
* NET 5156 = abc_8306_new_n1491
* NET 5158 = abc_8306_new_n1496
* NET 5160 = adrs[6]
* NET 5166 = abc_8306_new_n729
* NET 5171 = abc_8306_new_n371
* NET 5172 = abc_8306_new_n434
* NET 5173 = abc_8306_new_n370
* NET 5178 = abc_8306_new_n508
* NET 5181 = subckt_1571_sff1r_x4.sff_s
* NET 5185 = subckt_1571_sff1r_x4.sff_m
* NET 5188 = subckt_1571_sff1r_x4.ckr
* NET 5189 = subckt_1571_sff1r_x4.nckr
* NET 5207 = abc_8306_new_n317
* NET 5211 = abc_8306_new_n307
* NET 5212 = spare_buffer_170.q
* NET 5214 = abc_8306_new_n1625
* NET 5215 = abc_8306_new_n1626
* NET 5216 = data[3]
* NET 5218 = abc_8306_new_n1612
* NET 5220 = spare_buffer_166.q
* NET 5223 = spare_buffer_154.q
* NET 5225 = abc_8306_new_n323
* NET 5226 = abc_8306_new_n1224
* NET 5229 = abc_8306_auto_rtlil_cc_2608_muxgate_8127
* NET 5230 = abc_8306_new_n1579
* NET 5232 = spare_buffer_150.q
* NET 5233 = abc_8306_new_n1577
* NET 5234 = abc_8306_new_n1575
* NET 5235 = abc_8306_new_n1578
* NET 5238 = abc_8306_new_n1556
* NET 5239 = spare_buffer_90.q
* NET 5241 = abc_8306_new_n1530
* NET 5242 = abc_8306_new_n1540
* NET 5243 = abc_8306_new_n1539
* NET 5245 = spare_buffer_86.q
* NET 5247 = spare_buffer_74.q
* NET 5249 = abc_8306_new_n504
* NET 5251 = abc_8306_new_n1652
* NET 5252 = abc_8306_new_n536
* NET 5254 = spare_buffer_70.q
* NET 5256 = datao[6]
* NET 5267 = datao[0]
* NET 5268 = spare_buffer_169.q
* NET 5270 = m_clock_root_br_tr_br_0
* NET 5273 = abc_8306_new_n1282
* NET 5274 = data[2]
* NET 5275 = abc_8306_new_n1585
* NET 5278 = spare_buffer_165.q
* NET 5280 = m_clock_root_br_tr_0
* NET 5282 = abc_8306_new_n1417
* NET 5286 = abc_8306_new_n1637
* NET 5288 = spare_buffer_153.q
* NET 5291 = abc_8306_new_n1630
* NET 5294 = spare_buffer_149.q
* NET 5299 = abc_8306_new_n1507
* NET 5300 = abc_8306_new_n1512
* NET 5303 = spare_buffer_89.q
* NET 5306 = abc_8306_new_n730
* NET 5307 = abc_8306_new_n731
* NET 5310 = spare_buffer_85.q
* NET 5312 = m_clock_root_bl_tr_0
* NET 5317 = spare_buffer_73.q
* NET 5319 = spare_buffer_72.q
* NET 5325 = spare_buffer_69.q
* NET 5327 = m_clock_root_bl_tl_0
* NET 5329 = abc_8306_new_n242
* NET 5331 = abc_8306_auto_rtlil_cc_2608_muxgate_8067
* NET 5350 = adrs[10]
* NET 5351 = abc_8306_new_n1591
* NET 5352 = abc_8306_new_n1602
* NET 5353 = abc_8306_auto_rtlil_cc_2608_muxgate_8133
* NET 5355 = subckt_1609_sff1_x4.sff_s
* NET 5359 = subckt_1609_sff1_x4.sff_m
* NET 5361 = subckt_1609_sff1_x4.ckr
* NET 5362 = subckt_1609_sff1_x4.nckr
* NET 5364 = abc_8306_new_n1632
* NET 5365 = abc_8306_new_n1633
* NET 5366 = abc_8306_new_n1568
* NET 5369 = abc_8306_new_n1361
* NET 5371 = abc_8306_new_n290
* NET 5376 = abc_8306_new_n1360
* NET 5377 = abc_8306_new_n506
* NET 5378 = abc_8306_new_n503
* NET 5381 = abc_8306_new_n1472
* NET 5385 = abc_8306_new_n252
* NET 5386 = abc_8306_new_n485
* NET 5387 = abc_8306_new_n474
* NET 5393 = abc_8306_auto_rtlil_cc_2608_muxgate_8065
* NET 5411 = abc_8306_new_n1605
* NET 5413 = abc_8306_new_n1385
* NET 5417 = abc_8306_new_n1640
* NET 5418 = abc_8306_new_n1639
* NET 5420 = abc_8306_new_n1641
* NET 5421 = abc_8306_new_n1636
* NET 5423 = abc_8306_auto_rtlil_cc_2608_muxgate_8143
* NET 5425 = subckt_1599_sff1_x4.sff_s
* NET 5427 = subckt_1599_sff1_x4.sff_m
* NET 5429 = abc_8306_auto_rtlil_cc_2608_muxgate_8123
* NET 5432 = subckt_1599_sff1_x4.ckr
* NET 5433 = subckt_1599_sff1_x4.nckr
* NET 5434 = abc_8306_new_n1569
* NET 5435 = abc_8306_new_n322
* NET 5438 = abc_8306_new_n1513
* NET 5443 = subckt_1594_sff1_x4.sff_s
* NET 5444 = subckt_1594_sff1_x4.sff_m
* NET 5447 = subckt_1594_sff1_x4.ckr
* NET 5449 = m_clock_root_bl_tr_bl_0
* NET 5450 = subckt_1594_sff1_x4.nckr
* NET 5451 = abc_8306_new_n728
* NET 5454 = adrs[4]
* NET 5457 = abc_8306_new_n466
* NET 5459 = abc_8306_new_n1340
* NET 5460 = abc_8306_new_n1341
* NET 5461 = abc_8306_new_n1331
* NET 5466 = abc_8306_new_n479
* NET 5467 = abc_8306_new_n245
* NET 5470 = abc_8306_new_n241
* NET 5498 = abc_8306_new_n1603
* NET 5500 = abc_8306_new_n1606
* NET 5502 = abc_8306_new_n1607
* NET 5503 = abc_8306_new_n1426
* NET 5505 = abc_8306_new_n1392
* NET 5506 = abc_8306_new_n1383
* NET 5507 = abc_8306_new_n1424
* NET 5510 = subckt_1608_sff1_x4.sff_s
* NET 5513 = subckt_1608_sff1_x4.sff_m
* NET 5515 = abc_8306_auto_rtlil_cc_2608_muxgate_8141
* NET 5517 = subckt_1608_sff1_x4.ckr
* NET 5518 = m_clock_root_br_tl_bl_0
* NET 5519 = subckt_1608_sff1_x4.nckr
* NET 5520 = abc_8306_new_n1553
* NET 5521 = abc_8306_new_n1552
* NET 5523 = adrs[1]
* NET 5524 = subckt_1595_sff1_x4.sff_s
* NET 5528 = subckt_1595_sff1_x4.sff_m
* NET 5531 = m_clock_root_bl_tr_br_0
* NET 5532 = subckt_1595_sff1_x4.ckr
* NET 5533 = subckt_1595_sff1_x4.nckr
* NET 5534 = abc_8306_new_n1468
* NET 5535 = abc_8306_auto_rtlil_cc_2608_muxgate_8113
* NET 5536 = adrs[0]
* NET 5537 = abc_8306_new_n1190
* NET 5539 = abc_8306_new_n1191
* NET 5540 = datao[7]
* NET 5541 = abc_8306_new_n509
* NET 5544 = abc_8306_new_n384
* NET 5547 = subckt_1572_sff1r_x4.sff_s
* NET 5550 = subckt_1572_sff1r_x4.sff_m
* NET 5553 = subckt_1572_sff1r_x4.ckr
* NET 5554 = m_clock_root_bl_tl_bl_0
* NET 5555 = subckt_1572_sff1r_x4.nckr
* NET 5578 = subckt_1590_sff1_x4.sff_s
* NET 5581 = abc_8306_auto_rtlil_cc_2608_muxgate_8105
* NET 5582 = subckt_1590_sff1_x4.sff_m
* NET 5584 = m_clock_root_br_tr_bl_0
* NET 5585 = subckt_1590_sff1_x4.ckr
* NET 5587 = subckt_1590_sff1_x4.nckr
* NET 5589 = subckt_1592_sff1_x4.sff_s
* NET 5591 = subckt_1592_sff1_x4.sff_m
* NET 5594 = m_clock_root_br_tl_br_0
* NET 5595 = subckt_1592_sff1_x4.ckr
* NET 5597 = subckt_1592_sff1_x4.nckr
* NET 5600 = abc_8306_new_n1527
* NET 5604 = abc_8306_new_n1501
* NET 5606 = abc_8306_new_n294
* NET 5608 = abc_8306_new_n1073
* NET 5616 = abc_8306_new_n575
* NET 5617 = abc_8306_new_n578
* NET 5619 = abc_8306_new_n256
* NET 5620 = abc_8306_new_n469
* NET 5623 = sync
* NET 5625 = abc_8306_new_n1237
* NET 5626 = abc_8306_new_n1238
* NET 5653 = abc_8306_new_n302
* NET 5655 = abc_8306_new_n1405
* NET 5659 = abc_8306_new_n1414
* NET 5660 = abc_8306_new_n1407
* NET 5662 = abc_8306_new_n1364
* NET 5664 = abc_8306_new_n757
* NET 5667 = abc_8306_new_n1187
* NET 5669 = abc_8306_new_n1517
* NET 5670 = abc_8306_new_n1514
* NET 5671 = abc_8306_new_n1500
* NET 5675 = abc_8306_new_n1484
* NET 5676 = abc_8306_auto_rtlil_cc_2608_muxgate_8115
* NET 5677 = abc_8306_new_n1482
* NET 5678 = abc_8306_new_n1481
* NET 5679 = abc_8306_new_n1475
* NET 5681 = abc_8306_new_n911
* NET 5683 = abc_8306_new_n910
* NET 5685 = abc_8306_new_n1332
* NET 5688 = abc_8306_new_n1261
* NET 5690 = rdy_hfns_3
* NET 5691 = abc_8306_new_n468
* NET 5693 = abc_8306_new_n1229
* NET 5695 = abc_8306_new_n477
* NET 5706 = subckt_1587_sff1_x4.sff_m
* NET 5708 = abc_8306_new_n1448
* NET 5711 = abc_8306_new_n1528
* NET 5714 = subckt_1596_sff1_x4.sff_m
* NET 5716 = abc_8306_new_n1344
* NET 5718 = abc_8306_new_n380
* NET 5720 = abc_8306_new_n1227
* NET 5721 = subckt_1587_sff1_x4.sff_s
* NET 5723 = abc_8306_auto_rtlil_cc_2608_muxgate_8099
* NET 5725 = subckt_1587_sff1_x4.ckr
* NET 5726 = subckt_1587_sff1_x4.nckr
* NET 5727 = abc_8306_new_n1435
* NET 5728 = abc_8306_new_n1428
* NET 5729 = abc_8306_new_n1427
* NET 5734 = abc_8306_new_n1184
* NET 5735 = abc_8306_new_n1171
* NET 5738 = abc_8306_new_n1516
* NET 5739 = subckt_1596_sff1_x4.sff_s
* NET 5741 = abc_8306_auto_rtlil_cc_2608_muxgate_8117
* NET 5742 = subckt_1596_sff1_x4.ckr
* NET 5744 = subckt_1596_sff1_x4.nckr
* NET 5746 = adrs[5]
* NET 5751 = abc_8306_new_n1189
* NET 5757 = abc_8306_new_n1651
* NET 5792 = subckt_1591_sff1_x4.sff_s
* NET 5794 = subckt_1591_sff1_x4.sff_m
* NET 5797 = abc_8306_auto_rtlil_cc_2608_muxgate_8107
* NET 5799 = subckt_1591_sff1_x4.ckr
* NET 5800 = subckt_1591_sff1_x4.nckr
* NET 5801 = abc_8306_new_n1396
* NET 5803 = abc_8306_new_n1406
* NET 5804 = abc_8306_new_n1384
* NET 5805 = abc_8306_new_n1456
* NET 5806 = abc_8306_new_n1450
* NET 5807 = abc_8306_new_n1449
* NET 5809 = abc_8306_new_n1381
* NET 5810 = abc_8306_new_n912
* NET 5811 = abc_8306_new_n908
* NET 5812 = datao[1]
* NET 5813 = abc_8306_new_n1542
* NET 5815 = abc_8306_new_n1467
* NET 5816 = abc_8306_new_n1543
* NET 5817 = abc_8306_new_n312
* NET 5818 = abc_8306_new_n1471
* NET 5819 = abc_8306_new_n1474
* NET 5826 = abc_8306_new_n1470
* NET 5828 = abc_8306_new_n1485
* NET 5829 = abc_8306_new_n1498
* NET 5830 = abc_8306_new_n1497
* NET 5832 = abc_8306_new_n1259
* NET 5833 = adrs[7]
* NET 5834 = abc_8306_new_n1165
* NET 5835 = abc_8306_new_n1164
* NET 5837 = abc_8306_new_n1322
* NET 5840 = abc_8306_new_n465
* NET 5841 = ex_st_bit2_hfns_0
* NET 5842 = abc_8306_new_n473
* NET 5844 = abc_8306_new_n587
* NET 5846 = abc_8306_new_n1240
* NET 5848 = abc_8306_auto_rtlil_cc_2608_muxgate_8069
* NET 5860 = abc_8306_new_n276
* NET 5866 = subckt_1593_sff1_x4.sff_s
* NET 5870 = abc_8306_auto_rtlil_cc_2608_muxgate_8111
* NET 5871 = subckt_1593_sff1_x4.sff_m
* NET 5874 = subckt_1593_sff1_x4.nckr
* NET 5875 = subckt_1593_sff1_x4.ckr
* NET 5876 = abc_8306_new_n1328
* NET 5877 = abc_8306_new_n1348
* NET 5879 = abc_8306_new_n1437
* NET 5881 = abc_8306_auto_rtlil_cc_2608_muxgate_8109
* NET 5882 = dl[7]
* NET 5884 = abc_8306_new_n891
* NET 5885 = abc_8306_new_n905
* NET 5887 = dl[2]
* NET 5889 = abc_8306_new_n512
* NET 5891 = abc_8306_new_n1334
* NET 5895 = abc_8306_new_n1477
* NET 5897 = abc_8306_new_n727
* NET 5902 = abc_8306_new_n1327
* NET 5904 = abc_8306_new_n1343
* NET 5905 = abc_8306_new_n1342
* NET 5909 = abc_8306_new_n385
* NET 5912 = abc_8306_new_n478
* NET 5913 = abc_8306_new_n1225
* NET 5917 = abc_8306_new_n243
* NET 5944 = subckt_1588_sff1_x4.sff_s
* NET 5948 = subckt_1588_sff1_x4.sff_m
* NET 5950 = subckt_1588_sff1_x4.ckr
* NET 5951 = subckt_1588_sff1_x4.nckr
* NET 5952 = abc_8306_new_n1403
* NET 5953 = abc_8306_new_n1394
* NET 5954 = abc_8306_auto_rtlil_cc_2608_muxgate_8101
* NET 5955 = subckt_1586_sff1_x4.sff_s
* NET 5958 = subckt_1586_sff1_x4.sff_m
* NET 5960 = abc_8306_auto_rtlil_cc_2608_muxgate_8097
* NET 5963 = subckt_1586_sff1_x4.nckr
* NET 5964 = subckt_1586_sff1_x4.ckr
* NET 5966 = abc_8306_new_n1446
* NET 5967 = abc_8306_new_n1439
* NET 5969 = adrs[3]
* NET 5971 = subckt_1597_sff1_x4.sff_s
* NET 5974 = abc_8306_auto_rtlil_cc_2608_muxgate_8119
* NET 5976 = subckt_1597_sff1_x4.sff_m
* NET 5978 = subckt_1597_sff1_x4.nckr
* NET 5979 = subckt_1597_sff1_x4.ckr
* NET 5981 = abc_8306_new_n298
* NET 5982 = abc_8306_new_n590
* NET 5984 = abc_8306_new_n589
* NET 5985 = abc_8306_new_n588
* NET 5987 = abc_8306_new_n764
* NET 5988 = abc_8306_new_n760
* NET 5989 = abc_8306_new_n763
* NET 5991 = datao[5]
* NET 5992 = abc_8306_new_n1358
* NET 5994 = abc_8306_new_n461
* NET 6009 = abc_8306_new_n1617
* NET 6010 = abc_8306_new_n1419
* NET 6014 = abc_8306_new_n1421
* NET 6015 = abc_8306_new_n1423
* NET 6017 = abc_8306_new_n1416
* NET 6023 = abc_8306_new_n1363
* NET 6025 = dl[5]
* NET 6027 = abc_8306_new_n1140
* NET 6029 = abc_8306_new_n754
* NET 6030 = abc_8306_new_n713
* NET 6032 = abc_8306_new_n1672
* NET 6033 = abc_8306_new_n1667
* NET 6035 = dl[0]
* NET 6037 = abc_8306_new_n1670
* NET 6039 = abc_8306_new_n1074
* NET 6041 = abc_8306_new_n1075
* NET 6042 = abc_8306_new_n1072
* NET 6044 = abc_8306_new_n758
* NET 6046 = abc_8306_new_n1323
* NET 6047 = abc_8306_new_n1351
* NET 6048 = abc_8306_new_n1325
* NET 6056 = abc_8306_new_n1226
* NET 6058 = abc_8306_new_n1235
* NET 6061 = reg_762[2]
* NET 6094 = abc_8306_new_n1413
* NET 6096 = abc_8306_new_n1638
* NET 6099 = abc_8306_new_n1631
* NET 6102 = abc_8306_new_n1438
* NET 6107 = abc_8306_new_n1476
* NET 6111 = abc_8306_new_n1071
* NET 6112 = abc_8306_new_n1250
* NET 6114 = abc_8306_new_n1231
* NET 6115 = subckt_1589_sff1_x4.sff_s
* NET 6117 = subckt_1589_sff1_x4.sff_m
* NET 6119 = abc_8306_auto_rtlil_cc_2608_muxgate_8103
* NET 6120 = subckt_1589_sff1_x4.ckr
* NET 6121 = subckt_1589_sff1_x4.nckr
* NET 6124 = abc_8306_new_n1441
* NET 6125 = abc_8306_new_n364
* NET 6128 = abc_8306_new_n1049
* NET 6131 = abc_8306_new_n1143
* NET 6133 = ex_st_bit1_hfns_0
* NET 6135 = abc_8306_new_n244
* NET 6148 = spare_buffer_146.q
* NET 6150 = abc_8306_new_n1611
* NET 6154 = spare_buffer_142.q
* NET 6156 = abc_8306_new_n1362
* NET 6158 = abc_8306_new_n1395
* NET 6160 = abc_8306_new_n1451
* NET 6162 = abc_8306_new_n1455
* NET 6163 = spare_buffer_130.q
* NET 6165 = abc_8306_new_n1137
* NET 6166 = abc_8306_new_n1129
* NET 6168 = abc_8306_new_n941
* NET 6169 = abc_8306_new_n965
* NET 6172 = spare_buffer_126.q
* NET 6173 = dl[6]
* NET 6175 = dl[4]
* NET 6177 = spare_buffer_66.q
* NET 6180 = abc_8306_new_n1469
* NET 6181 = abc_8306_new_n585
* NET 6183 = spare_buffer_62.q
* NET 6185 = abc_8306_new_n909
* NET 6187 = adrs[2]
* NET 6191 = spare_buffer_50.q
* NET 6193 = abc_8306_new_n1350
* NET 6194 = abc_8306_new_n1262
* NET 6195 = abc_8306_new_n1349
* NET 6199 = spare_buffer_46.q
* NET 6202 = abc_8306_new_n1309
* NET 6222 = spare_buffer_145.q
* NET 6226 = abc_8306_new_n1422
* NET 6229 = spare_buffer_141.q
* NET 6231 = m_clock_root_br_br_tl_0
* NET 6234 = abc_8306_new_n1453
* NET 6237 = spare_buffer_129.q
* NET 6241 = abc_8306_new_n1702
* NET 6242 = abc_8306_new_n1687
* NET 6243 = spare_buffer_125.q
* NET 6246 = abc_8306_new_n1707
* NET 6247 = abc_8306_new_n1682
* NET 6249 = spare_buffer_65.q
* NET 6253 = abc_8306_new_n581
* NET 6254 = spare_buffer_61.q
* NET 6256 = spare_buffer_60.q
* NET 6259 = abc_8306_new_n952
* NET 6261 = spare_buffer_49.q
* NET 6263 = spare_buffer_48.q
* NET 6266 = ex_st[0]
* NET 6267 = abc_8306_new_n464
* NET 6268 = spare_buffer_45.q
* NET 6271 = abc_8306_new_n1307
* NET 6272 = abc_8306_new_n1311
* NET 6291 = abc_8306_new_n1412
* NET 6293 = abc_8306_new_n1408
* NET 6296 = subckt_1631_sff1_x4.sff_s
* NET 6300 = subckt_1631_sff1_x4.sff_m
* NET 6302 = m_clock_root_br_bl_tr_0
* NET 6303 = subckt_1631_sff1_x4.ckr
* NET 6305 = subckt_1631_sff1_x4.nckr
* NET 6306 = abc_8306_new_n1709
* NET 6309 = abc_8306_new_n1712
* NET 6310 = abc_8306_new_n1710
* NET 6314 = abc_8306_new_n928
* NET 6315 = abc_8306_new_n1666
* NET 6316 = abc_8306_new_n918
* NET 6318 = abc_8306_new_n1695
* NET 6322 = abc_8306_new_n1671
* NET 6323 = abc_8306_new_n264
* NET 6325 = abc_8306_new_n1050
* NET 6326 = abc_8306_new_n1051
* NET 6328 = abc_8306_new_n1163
* NET 6332 = abc_8306_new_n463
* NET 6333 = rdy_hfns_1
* NET 6336 = abc_8306_new_n1335
* NET 6337 = abc_8306_new_n535
* NET 6338 = abc_8306_new_n586
* NET 6339 = abc_8306_new_n1288
* NET 6340 = abc_8306_new_n1278
* NET 6341 = abc_8306_new_n1312
* NET 6342 = abc_8306_new_n1270
* NET 6344 = abc_8306_new_n327
* NET 6372 = abc_8306_new_n1411
* NET 6375 = abc_8306_new_n1418
* NET 6378 = abc_8306_new_n1434
* NET 6380 = abc_8306_new_n1452
* NET 6382 = abc_8306_new_n1445
* NET 6384 = abc_8306_new_n1716
* NET 6386 = abc_8306_new_n1524
* NET 6388 = dl[3]
* NET 6389 = abc_8306_new_n1689
* NET 6391 = abc_8306_new_n1669
* NET 6392 = dl[1]
* NET 6393 = abc_8306_new_n1359
* NET 6394 = abc_8306_new_n1333
* NET 6397 = abc_8306_new_n811
* NET 6399 = abc_8306_new_n809
* NET 6400 = abc_8306_new_n810
* NET 6402 = abc_8306_new_n1048
* NET 6405 = abc_8306_new_n1338
* NET 6406 = abc_8306_new_n1377
* NET 6407 = abc_8306_new_n362
* NET 6408 = abc_8306_new_n352
* NET 6409 = wt
* NET 6410 = nmi
* NET 6432 = ry[5]
* NET 6434 = subckt_1663_sff1_x4.sff_s
* NET 6436 = subckt_1663_sff1_x4.sff_m
* NET 6439 = abc_8306_auto_rtlil_cc_2608_muxgate_8283
* NET 6441 = subckt_1663_sff1_x4.ckr
* NET 6442 = subckt_1663_sff1_x4.nckr
* NET 6443 = abc_8306_new_n271
* NET 6444 = abc_8306_new_n1597
* NET 6451 = abc_8306_new_n1574
* NET 6456 = subckt_1627_sff1_x4.sff_s
* NET 6458 = subckt_1627_sff1_x4.sff_m
* NET 6462 = subckt_1627_sff1_x4.ckr
* NET 6463 = subckt_1627_sff1_x4.nckr
* NET 6464 = abc_8306_new_n1674
* NET 6466 = abc_8306_auto_rtlil_cc_2608_muxgate_8179
* NET 6469 = abc_8306_new_n1006
* NET 6471 = abc_8306_new_n1162
* NET 6473 = abc_8306_new_n951
* NET 6474 = abc_8306_new_n363
* NET 6476 = datao[4]
* NET 6477 = abc_8306_new_n1330
* NET 6482 = subckt_1667_sff1r_x4.sff_s
* NET 6486 = subckt_1667_sff1r_x4.sff_m
* NET 6489 = subckt_1667_sff1r_x4.ckr
* NET 6490 = subckt_1667_sff1r_x4.nckr
* NET 6491 = nm1
* NET 6518 = abc_8306_new_n1399
* NET 6519 = abc_8306_new_n1409
* NET 6521 = abc_8306_new_n1454
* NET 6523 = abc_8306_new_n1440
* NET 6528 = m_clock_root_br_bl_tl_0
* NET 6529 = abc_8306_new_n1492
* NET 6531 = abc_8306_new_n808
* NET 6532 = abc_8306_new_n1005
* NET 6533 = abc_8306_new_n386
* NET 6534 = abc_8306_new_n1222
* NET 6535 = abc_8306_new_n1234
* NET 6538 = abc_8306_new_n1230
* NET 6539 = adrs[13]
* NET 6540 = subckt_1607_sff1_x4.sff_s
* NET 6542 = subckt_1607_sff1_x4.sff_m
* NET 6544 = subckt_1607_sff1_x4.ckr
* NET 6545 = subckt_1607_sff1_x4.nckr
* NET 6549 = abc_8306_auto_rtlil_cc_2608_muxgate_8139
* NET 6553 = abc_8306_new_n1442
* NET 6555 = subckt_1632_sff1_x4.sff_s
* NET 6556 = subckt_1632_sff1_x4.ckr
* NET 6557 = subckt_1632_sff1_x4.nckr
* NET 6559 = subckt_1632_sff1_x4.sff_m
* NET 6561 = abc_8306_auto_rtlil_cc_2608_muxgate_8189
* NET 6562 = abc_8306_new_n1683
* NET 6565 = abc_8306_new_n583
* NET 6566 = abc_8306_new_n582
* NET 6568 = abc_8306_new_n1004
* NET 6569 = abc_8306_new_n1003
* NET 6570 = abc_8306_new_n833
* NET 6572 = abc_8306_new_n834
* NET 6576 = abc_8306_new_n1233
* NET 6590 = subckt_1661_sff1_x4.sff_m
* NET 6592 = subckt_1661_sff1_x4.ckr
* NET 6593 = abc_8306_new_n1700
* NET 6594 = abc_8306_auto_rtlil_cc_2608_muxgate_8187
* NET 6596 = abc_8306_new_n1680
* NET 6598 = abc_8306_new_n1685
* NET 6599 = abc_8306_new_n1352
* NET 6600 = abc_8306_new_n1258
* NET 6606 = subckt_1580_sff1r_x4.sff_m
* NET 6608 = abc_8306_auto_rtlil_cc_2608_muxgate_8085
* NET 6610 = subckt_1580_sff1r_x4.ckr
* NET 6611 = m_clock_root_bl_bl_tl_0
* NET 6612 = subckt_1580_sff1r_x4.nckr
* NET 6613 = abc_8306_auto_rtlil_cc_2608_muxgate_8291
* NET 6614 = abc_8306_new_n1765
* NET 6616 = subckt_1661_sff1_x4.sff_s
* NET 6617 = ry[3]
* NET 6619 = subckt_1661_sff1_x4.nckr
* NET 6620 = abc_8306_auto_rtlil_cc_2608_muxgate_8279
* NET 6622 = m_clock_root_br_br_tr_0
* NET 6625 = abc_8306_new_n1432
* NET 6628 = debug[15]
* NET 6629 = abc_8306_new_n285
* NET 6631 = abc_8306_new_n1390
* NET 6632 = abc_8306_new_n1692
* NET 6633 = abc_8306_new_n1690
* NET 6637 = abc_8306_new_n1522
* NET 6641 = abc_8306_new_n1681
* NET 6644 = abc_8306_new_n835
* NET 6646 = abc_8306_new_n836
* NET 6648 = abc_8306_new_n1508
* NET 6651 = subckt_1580_sff1r_x4.sff_s
* NET 6652 = int_req
* NET 6672 = abc_8306_new_n1624
* NET 6676 = debug[14]
* NET 6678 = abc_8306_new_n1444
* NET 6681 = abc_8306_new_n1714
* NET 6682 = abc_8306_new_n1705
* NET 6683 = abc_8306_new_n1703
* NET 6685 = subckt_1626_sff1_x4.sff_s
* NET 6688 = subckt_1626_sff1_x4.sff_m
* NET 6690 = abc_8306_auto_rtlil_cc_2608_muxgate_8177
* NET 6693 = m_clock_root_bl_br_tr_0
* NET 6694 = subckt_1626_sff1_x4.nckr
* NET 6695 = subckt_1626_sff1_x4.ckr
* NET 6696 = abc_8306_new_n1675
* NET 6697 = abc_8306_new_n1678
* NET 6698 = abc_8306_new_n1676
* NET 6700 = abc_8306_new_n953
* NET 6703 = abc_8306_new_n954
* NET 6704 = abc_8306_new_n1145
* NET 6705 = abc_8306_new_n1144
* NET 6707 = abc_8306_new_n1019
* NET 6708 = abc_8306_new_n762
* NET 6710 = abc_8306_new_n395
* NET 6713 = abc_8306_new_n1317
* NET 6714 = abc_8306_new_n366
* NET 6726 = abc_8306_new_n1410
* NET 6731 = abc_8306_new_n1430
* NET 6732 = abc_8306_new_n279
* NET 6733 = abc_8306_new_n282
* NET 6736 = abc_8306_new_n1443
* NET 6739 = m_clock_root_br_0
* NET 6741 = abc_8306_new_n1688
* NET 6745 = subckt_1628_sff1_x4.sff_s
* NET 6749 = subckt_1628_sff1_x4.sff_m
* NET 6750 = abc_8306_auto_rtlil_cc_2608_muxgate_8181
* NET 6752 = subckt_1628_sff1_x4.ckr
* NET 6753 = subckt_1628_sff1_x4.nckr
* NET 6757 = abc_8306_new_n1047
* NET 6761 = abc_8306_new_n968
* NET 6762 = datao[3]
* NET 6764 = abc_8306_new_n1142
* NET 6768 = abc_8306_new_n392
* NET 6770 = abc_8306_new_n262
* NET 6771 = m_clock_root_bl_0
* NET 6773 = abc_8306_new_n1228
* NET 6804 = rx[5]
* NET 6806 = subckt_1655_sff1_x4.sff_s
* NET 6810 = subckt_1655_sff1_x4.sff_m
* NET 6811 = abc_8306_auto_rtlil_cc_2608_muxgate_8267
* NET 6813 = subckt_1655_sff1_x4.ckr
* NET 6814 = subckt_1655_sff1_x4.nckr
* NET 6817 = abc_8306_new_n1433
* NET 6819 = abc_8306_new_n1431
* NET 6822 = subckt_1629_sff1_x4.sff_s
* NET 6825 = abc_8306_auto_rtlil_cc_2608_muxgate_8183
* NET 6827 = subckt_1629_sff1_x4.sff_m
* NET 6829 = subckt_1629_sff1_x4.ckr
* NET 6830 = subckt_1629_sff1_x4.nckr
* NET 6831 = abc_8306_new_n1708
* NET 6832 = abc_8306_new_n1561
* NET 6836 = abc_8306_new_n1696
* NET 6837 = abc_8306_new_n1694
* NET 6839 = abc_8306_new_n1494
* NET 6840 = abc_8306_new_n832
* NET 6841 = abc_8306_new_n950
* NET 6843 = abc_8306_new_n1329
* NET 6845 = abc_8306_new_n261
* NET 6846 = abc_8306_new_n375
* NET 6848 = abc_8306_new_n1354
* NET 6849 = abc_8306_new_n1220
* NET 6851 = abc_8306_new_n1764
* NET 6852 = abc_8306_new_n1218
* NET 6869 = abc_8306_new_n1420
* NET 6876 = abc_8306_new_n1719
* NET 6878 = abc_8306_new_n1717
* NET 6882 = abc_8306_new_n1701
* NET 6885 = abc_8306_new_n1521
* NET 6886 = abc_8306_new_n1560
* NET 6888 = abc_8306_new_n1535
* NET 6892 = abc_8306_new_n1698
* NET 6893 = abc_8306_new_n1665
* NET 6894 = abc_8306_new_n1015
* NET 6897 = abc_8306_new_n807
* NET 6899 = abc_8306_new_n1141
* NET 6901 = abc_8306_new_n1023
* NET 6902 = abc_8306_new_n1022
* NET 6906 = abc_8306_new_n388
* NET 6907 = abc_8306_new_n382
* NET 6910 = abc_8306_new_n1221
* NET 6912 = abc_8306_new_n1219
* NET 6914 = abc_8306_new_n1493
* NET 6917 = abc_8306_new_n369
* NET 6940 = abc_8306_new_n1402
* NET 6942 = abc_8306_new_n1429
* NET 6944 = abc_8306_new_n1584
* NET 6947 = abc_8306_new_n1715
* NET 6948 = abc_8306_new_n1691
* NET 6954 = abc_8306_new_n1002
* NET 6955 = abc_8306_new_n1188
* NET 6957 = abc_8306_new_n1510
* NET 6965 = debug[13]
* NET 6967 = abc_8306_new_n1668
* NET 6968 = abc_8306_new_n1357
* NET 6969 = abc_8306_new_n1520
* NET 6971 = subckt_1630_sff1_x4.sff_s
* NET 6973 = subckt_1630_sff1_x4.sff_m
* NET 6974 = subckt_1630_sff1_x4.nckr
* NET 6976 = abc_8306_auto_rtlil_cc_2608_muxgate_8185
* NET 6977 = subckt_1630_sff1_x4.ckr
* NET 6979 = abc_8306_new_n577
* NET 6980 = abc_8306_new_n576
* NET 6981 = abc_8306_new_n1223
* NET 6982 = subckt_1582_sff1r_x4.sff_s
* NET 6983 = subckt_1582_sff1r_x4.nckr
* NET 6985 = subckt_1582_sff1r_x4.sff_m
* NET 6987 = subckt_1582_sff1r_x4.ckr
* NET 6988 = abc_8306_auto_rtlil_cc_2608_muxgate_8089
* NET 6990 = abc_8306_new_n1308
* NET 6991 = do_brk
* NET 6992 = abc_8306_new_n324
* NET 7010 = abc_8306_new_n1604
* NET 7011 = abc_8306_new_n1401
* NET 7016 = abc_8306_new_n1379
* NET 7018 = abc_8306_new_n1548
* NET 7024 = abc_8306_new_n1519
* NET 7027 = abc_8306_new_n1506
* NET 7031 = abc_8306_new_n1490
* NET 7032 = abc_8306_new_n1355
* NET 7033 = abc_8306_new_n1353
* NET 7034 = abc_8306_new_n1376
* NET 7039 = abc_8306_new_n1017
* NET 7042 = ex_st_bit2_hfns_1
* NET 7044 = abc_8306_new_n387
* NET 7045 = abc_8306_new_n1316
* NET 7049 = abc_8306_new_n1216
* NET 7074 = abc_8306_new_n1386
* NET 7075 = abc_8306_new_n1400
* NET 7078 = abc_8306_new_n1398
* NET 7082 = subckt_1633_sff1_x4.sff_s
* NET 7084 = abc_8306_auto_rtlil_cc_2608_muxgate_8191
* NET 7085 = subckt_1633_sff1_x4.sff_m
* NET 7088 = subckt_1633_sff1_x4.nckr
* NET 7089 = subckt_1633_sff1_x4.ckr
* NET 7092 = abc_8306_new_n1518
* NET 7094 = abc_8306_new_n272
* NET 7095 = abc_8306_new_n1366
* NET 7098 = abc_8306_new_n1697
* NET 7099 = abc_8306_new_n1505
* NET 7101 = abc_8306_new_n1489
* NET 7103 = abc_8306_new_n970
* NET 7104 = abc_8306_new_n972
* NET 7105 = abc_8306_new_n971
* NET 7107 = abc_8306_new_n931
* NET 7108 = ex_st[3]
* NET 7109 = abc_8306_new_n376
* NET 7110 = abc_8306_new_n394
* NET 7111 = abc_8306_new_n326
* NET 7113 = abc_8306_new_n325
* NET 7114 = rdy_hfns_0
* NET 7123 = datao[2]
* NET 7124 = spare_buffer_138.q
* NET 7126 = spare_buffer_134.q
* NET 7129 = abc_8306_new_n1388
* NET 7133 = spare_buffer_122.q
* NET 7137 = abc_8306_new_n1571
* NET 7141 = spare_buffer_118.q
* NET 7144 = abc_8306_new_n1533
* NET 7147 = spare_buffer_58.q
* NET 7149 = abc_8306_new_n1677
* NET 7151 = abc_8306_new_n1488
* NET 7154 = spare_buffer_54.q
* NET 7156 = abc_8306_new_n969
* NET 7160 = spare_buffer_42.q
* NET 7162 = rdy_hfns_2
* NET 7163 = abc_8306_new_n1232
* NET 7164 = abc_8306_new_n476
* NET 7168 = abc_8306_new_n1217
* NET 7170 = spare_buffer_38.q
* NET 7173 = abc_8306_new_n275
* NET 7174 = abc_8306_new_n1315
* NET 7187 = spare_buffer_137.q
* NET 7189 = m_clock_root_br_br_br_0
* NET 7191 = spare_buffer_133.q
* NET 7193 = spare_buffer_132.q
* NET 7194 = m_clock_root_br_br_0
* NET 7196 = abc_8306_new_n268
* NET 7197 = spare_buffer_121.q
* NET 7199 = m_clock_root_br_bl_br_0
* NET 7205 = spare_buffer_117.q
* NET 7208 = m_clock_root_br_bl_bl_0
* NET 7210 = abc_8306_new_n1559
* NET 7212 = abc_8306_new_n1711
* NET 7213 = spare_buffer_57.q
* NET 7215 = m_clock_root_bl_br_br_0
* NET 7218 = abc_8306_new_n1684
* NET 7219 = abc_8306_new_n1504
* NET 7222 = spare_buffer_53.q
* NET 7224 = m_clock_root_bl_br_0
* NET 7225 = m_clock_root_bl_br_bl_0
* NET 7227 = abc_8306_new_n393
* NET 7228 = abc_8306_new_n390
* NET 7230 = spare_buffer_41.q
* NET 7232 = spare_buffer_40.q
* NET 7234 = abc_8306_new_n1021
* NET 7235 = ift_run
* NET 7236 = abc_8306_new_n1215
* NET 7238 = spare_buffer_37.q
* NET 7242 = abc_8306_new_n1310
* NET 7243 = abc_8306_new_n1319
* NET 7255 = abc_8306_new_n1397
* NET 7261 = abc_8306_new_n1378
* NET 7263 = abc_8306_new_n1380
* NET 7264 = abc_8306_new_n1718
* NET 7267 = abc_8306_new_n1573
* NET 7270 = abc_8306_new_n1557
* NET 7274 = abc_8306_new_n1532
* NET 7278 = abc_8306_new_n1534
* NET 7280 = abc_8306_new_n1375_hfns_1
* NET 7283 = abc_8306_new_n1339
* NET 7286 = abc_8306_new_n383
* NET 7287 = abc_8306_new_n254
* NET 7289 = abc_8306_new_n1509
* NET 7307 = abc_8306_new_n1374
* NET 7309 = abc_8306_new_n1572
* NET 7311 = abc_8306_new_n1547
* NET 7313 = abc_8306_new_n1558
* NET 7315 = abc_8306_new_n1486
* NET 7317 = abc_8306_new_n1487
* NET 7320 = abc_8306_new_n1018
* NET 7334 = abc_8306_new_n377
* NET 7335 = debug[12]
* NET 7337 = subckt_1584_sff1r_x4.sff_s
* NET 7339 = subckt_1584_sff1r_x4.sff_m
* NET 7341 = subckt_1584_sff1r_x4.ckr
* NET 7342 = subckt_1584_sff1r_x4.nckr
* NET 7343 = abc_8306_auto_rtlil_cc_2608_muxgate_8093
* NET 7353 = abc_8306_new_n389
* NET 7354 = abc_8306_new_n391
* NET 7356 = abc_8306_new_n1020
* NET 7357 = abc_8306_new_n1389
* NET 7358 = abc_8306_new_n1391
* NET 7366 = abc_8306_new_n1545
* NET 7369 = abc_8306_new_n277
* NET 7372 = abc_8306_new_n1531
* NET 7377 = abc_8306_new_n1502
* NET 7379 = abc_8306_new_n1339_hfns_0
* NET 7381 = abc_8306_new_n1375
* NET 7383 = abc_8306_new_n368
* NET 7384 = abc_8306_new_n365
* NET 7387 = do_nmi
* NET 7388 = reg_762[0]
* NET 7390 = reg_762[1]
* NET 7391 = abc_8306_new_n367
* NET 7411 = abc_8306_new_n1373
* NET 7413 = abc_8306_new_n1371
* NET 7416 = abc_8306_new_n1570
* NET 7418 = abc_8306_new_n1370
* NET 7419 = abc_8306_new_n1546
* NET 7420 = abc_8306_new_n1356
* NET 7422 = abc_8306_new_n1704
* NET 7424 = abc_8306_new_n283
* NET 7427 = abc_8306_new_n1339_hfns_2
* NET 7428 = abc_8306_new_n1339_hfns_1
* NET 7430 = abc_8306_new_n932
* NET 7431 = abc_8306_new_n935
* NET 7432 = abc_8306_new_n934
* NET 7433 = abc_8306_new_n933
* NET 7436 = subckt_1583_sff1r_x4.sff_s
* NET 7439 = subckt_1583_sff1r_x4.sff_m
* NET 7440 = abc_8306_auto_rtlil_cc_2608_muxgate_8091
* NET 7443 = subckt_1583_sff1r_x4.ckr
* NET 7444 = subckt_1583_sff1r_x4.nckr
* NET 7451 = vdd
* NET 7452 = debug[11]
* NET 7453 = debug[10]
* NET 7454 = debug[9]
* NET 7455 = abc_8306_new_n266
* NET 7458 = abc_8306_new_n1387
* NET 7460 = abc_8306_new_n1372
* NET 7462 = debug[8]
* NET 7463 = abc_8306_new_n263
* NET 7464 = debug[7]
* NET 7465 = abc_8306_new_n286
* NET 7466 = debug[6]
* NET 7470 = abc_8306_new_n1544
* NET 7471 = abc_8306_new_n1368
* NET 7473 = abc_8306_new_n280
* NET 7474 = abc_8306_new_n1369
* NET 7475 = debug[5]
* NET 7477 = abc_8306_new_n1367
* NET 7480 = debug[4]
* NET 7481 = debug[3]
* NET 7484 = abc_8306_new_n1503
* NET 7486 = abc_8306_new_n1365
* NET 7488 = abc_8306_new_n269
* NET 7489 = debug[2]
* NET 7490 = abc_8306_new_n1375_hfns_2
* NET 7491 = abc_8306_new_n1375_hfns_0
* NET 7493 = debug[1]
* NET 7494 = debug[0]
* NET 7495 = adrs[15]
* NET 7496 = do_res
* NET 7499 = subckt_1581_sff1r_x4.sff_s
* NET 7500 = p_reset_hfns_0
* NET 7504 = subckt_1581_sff1r_x4.sff_m
* NET 7505 = abc_8306_auto_rtlil_cc_2608_muxgate_8087
* NET 7508 = m_clock_root_bl_bl_bl_0
* NET 7509 = subckt_1581_sff1r_x4.nckr
* NET 7510 = subckt_1581_sff1r_x4.ckr
* NET 7511 = adrs[14]
* NET 7512 = do_irq
* NET 7513 = abc_8306_new_n274
* NET 7514 = vss
Mtr_16378 7451 7240 7171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16377 7170 7171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16376 7451 7171 7170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16375 7451 7171 7170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16374 7170 7171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16373 1169 1449 4446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16372 1170 1168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16371 7451 1170 1169 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16370 3067 2922 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16369 3067 2645 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16368 7451 2412 3067 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16367 356 1021 357 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_16366 355 1023 356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_16365 7451 1022 355 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_16364 1020 357 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16363 5563 6316 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16362 5671 6314 5563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16361 7451 5815 5671 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16360 7451 7240 7239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16359 7238 7239 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16358 7451 7239 7238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16357 7451 7239 7238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16356 7238 7239 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16355 7451 7240 7241 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16354 7508 7241 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16353 7451 7241 7508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16352 7451 7241 7508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16351 7508 7241 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16350 7451 6771 4776 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16349 5312 4776 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16348 7451 4776 5312 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16347 7451 4776 5312 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16346 5312 4776 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16345 6279 6316 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16344 6596 6314 6279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16343 7451 6315 6596 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16342 3107 3581 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16341 7451 3107 3105 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16340 3106 3324 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16339 7451 3106 3103 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16338 3103 3105 3104 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16337 3104 3107 3102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16336 3099 4424 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_16335 7451 3100 4424 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16334 4424 3100 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16333 3102 3101 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16332 3101 3104 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16331 7451 5100 3101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16330 3100 5100 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16329 3100 3105 3099 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_16328 3101 3107 3100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_16327 7451 6771 4788 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16326 5327 4788 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16325 7451 4788 5327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16324 7451 4788 5327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16323 5327 4788 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16322 7451 6771 6756 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16321 7224 6756 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16320 7451 6756 7224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16319 7451 6756 7224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16318 7224 6756 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16317 7451 6771 6772 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16316 7240 6772 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16315 7451 6772 7240 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16314 7451 6772 7240 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16313 7240 6772 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16312 1654 1832 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16311 7451 4588 1654 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16310 1653 1654 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16309 6908 7044 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16308 7451 6907 6908 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16307 6906 6908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16306 2660 3149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16305 2661 4695 2660 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16304 7451 2856 2661 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16303 7385 7391 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16302 7451 7384 7385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16301 7383 7385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16300 7451 5752 1739 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16299 2712 1739 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16298 7451 1739 2712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16297 7451 1739 2712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16296 2712 1739 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16295 7451 5752 1762 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16294 2746 1762 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16293 7451 1762 2746 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16292 7451 1762 2746 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16291 2746 1762 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16290 7451 1040 713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16289 713 1041 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16288 713 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16287 7451 4589 713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16286 832 713 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16285 71 72 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16284 67 73 66 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16283 7451 4104 67 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16282 73 74 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_16281 7451 368 74 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_16280 7451 4103 72 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16279 69 73 71 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16278 70 74 69 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16277 7451 68 70 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16276 68 69 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16275 66 74 68 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16274 7451 66 4104 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16273 4104 66 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16272 7451 5171 4935 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16271 4935 5172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16270 4935 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16269 7451 7042 4935 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16268 6566 4935 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16267 7451 4161 727 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16266 727 1168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16265 7451 4376 727 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16264 1292 727 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16263 5666 5734 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16262 5667 5735 5666 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16261 7451 6125 5667 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16260 6314 3562 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16259 7451 3563 6314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16258 3804 3487 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16257 7451 3409 3804 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16256 2293 2292 2276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16255 2276 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16254 7451 2392 2276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16253 2652 2293 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16252 2275 2583 2293 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16251 2276 3549 2275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16250 6385 6384 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16249 7451 6386 6385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16248 6878 6385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16247 4686 5215 4702 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16246 4703 4701 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16245 7451 4703 4686 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16244 4978 4975 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16243 4978 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16242 7451 5826 4978 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16241 638 3546 639 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16240 639 2576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16239 7451 1851 639 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16238 1679 638 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16237 637 3549 638 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16236 639 3545 637 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16235 5260 5417 5420 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16234 5287 5286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16233 7451 5287 5260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16232 4847 4642 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16231 4847 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16230 7451 5826 4847 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16229 3343 5138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16228 3343 3655 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16227 7451 3170 3343 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16226 4240 4841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16225 4257 4413 4240 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16224 4239 4411 4257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16223 7451 4255 4239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16222 4254 4257 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16221 2404 2416 2405 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16220 2405 2418 2419 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16219 2419 2789 2405 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16218 2404 2504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16217 7451 2424 2404 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16216 2405 2502 2404 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16215 2648 2419 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16214 7326 7379 7310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16213 7310 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16212 7451 7464 7326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16211 7309 7326 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16210 2316 2676 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16209 7451 2956 2316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16208 2315 2316 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16207 1985 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16206 2228 2929 1985 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16205 7451 6175 2228 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16204 1818 2023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16203 7451 2288 1818 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16202 1821 1818 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16201 2959 2988 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16200 7451 2958 2959 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16199 3030 2959 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16198 7451 5459 5463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16197 5463 5460 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16196 5463 6405 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16195 7451 5461 5463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16194 5905 5463 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16193 7451 5891 5890 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16192 5890 5992 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16191 5890 5902 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16190 7451 5889 5890 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16189 6156 5890 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16188 2549 2552 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16187 2545 2551 2546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16186 7451 7108 2545 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16185 2551 2554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_16184 7451 2553 2554 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_16183 7451 2752 2552 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16182 2550 2551 2549 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16181 2548 2554 2550 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16180 7451 2547 2548 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16179 2547 2550 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16178 2546 2554 2547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16177 7451 2546 7108 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16176 7108 2546 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16175 4678 5691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16174 7451 7108 4678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16173 4679 4678 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16172 7237 7387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16171 7236 7512 7237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16170 7451 7235 7236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16169 7037 7101 7002 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16168 7002 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16167 7451 7034 7002 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16166 7031 7037 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16165 7001 7032 7037 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16164 7002 7317 7001 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16163 7451 6518 6292 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16162 6291 7452 6274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16161 6274 6518 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16160 6274 6292 6291 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16159 7451 6289 6274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16158 6289 7452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16157 5261 6030 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16156 5534 6029 5261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16155 7451 5815 5534 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16154 7451 1872 1873 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16153 1873 1871 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16152 7451 2798 1873 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16151 2018 1873 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16150 1498 1834 1463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16149 1463 1620 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16148 7451 1619 1463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16147 1496 1498 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16146 1462 3425 1498 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16145 1463 1631 1462 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16144 7451 5842 3928 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16143 3928 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16142 7451 5690 3928 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16141 3927 3928 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16140 7451 1435 904 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16139 904 1768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16138 903 902 904 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16137 901 899 903 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16136 904 900 901 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16135 4752 4837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16134 7451 6009 4752 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16133 7451 2748 2734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16132 2734 2741 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16131 2734 5093 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16130 7451 4732 2734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16129 2733 2734 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16128 7451 6565 5086 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16127 5086 6566 5085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16126 4966 4758 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16125 7451 4195 4966 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16124 4754 5218 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16123 7451 6150 4754 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16122 652 960 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16121 777 832 652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16120 7451 2592 777 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16119 1340 1605 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16118 7451 1426 1340 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16117 6342 5623 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16116 7451 6333 6342 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16115 2973 2971 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16114 2973 2972 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16113 7451 3259 2973 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16112 3415 6030 3713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16111 3416 3957 3415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16110 7451 3958 3416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16109 4827 5097 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16108 7451 4829 4827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16107 7451 181 179 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16106 563 509 182 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16105 182 181 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16104 182 179 563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16103 7451 180 182 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16102 180 509 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16101 2931 3135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16100 7451 3500 2931 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16099 5267 5987 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16098 7451 5664 5267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16097 924 2139 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16096 939 3545 924 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16095 7451 1688 939 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16094 6479 6843 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16093 7451 6907 6479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16092 6477 6479 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16091 6158 7453 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16090 6158 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16089 7451 6968 6158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16088 7451 894 502 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16087 3409 691 504 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16086 504 894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16085 504 502 3409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16084 7451 503 504 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16083 503 691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16082 1414 3545 1415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16081 1415 2095 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16080 7451 1688 1414 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16079 1413 1414 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16078 7451 5913 5758 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16077 5758 5844 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16076 7451 6267 5758 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16075 5757 5758 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16074 2925 2102 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16073 2925 2318 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16072 7451 2171 2925 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16071 7451 4773 2925 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16070 4674 2881 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16069 4674 2880 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16068 7451 4446 4674 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16067 4766 5275 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16066 4848 5273 4766 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16065 7451 5043 4848 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16064 1820 1823 1822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16063 1822 1821 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16062 7451 2154 1820 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16061 1819 1820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16060 3574 3571 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16059 7451 3574 3572 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16058 3573 3568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16057 7451 3573 3569 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16056 3569 3572 3570 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16055 3570 3574 3567 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16054 3564 4991 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_16053 7451 3565 4991 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16052 4991 3565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16051 3567 3566 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16050 3566 3570 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16049 7451 7500 3566 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16048 3565 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16047 3565 3572 3564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_16046 3566 3574 3565 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_16045 2413 4695 2403 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16044 2403 3129 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16043 7451 3128 2413 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16042 2412 2413 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_16041 5674 5743 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16040 5672 5742 5739 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16039 7451 6187 5672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16038 5742 5744 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_16037 7451 6693 5744 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_16036 7451 5741 5743 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16035 5714 5742 5674 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16034 5673 5744 5714 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16033 7451 5713 5673 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16032 5713 5714 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16031 5739 5744 5713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_16030 7451 5739 6187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16029 6187 5739 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16028 187 2016 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16027 7451 3546 187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16026 186 187 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16025 7451 1029 689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16024 689 1145 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16023 7451 1809 689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16022 1021 689 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16021 1436 2174 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16020 1435 1837 1436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16019 7451 6333 1435 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16018 1386 1385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16017 7451 1384 1386 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16016 2033 1386 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16015 7451 7095 7022 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16014 7024 7481 6998 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16013 6998 7095 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16012 6998 7022 7024 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16011 7451 7023 6998 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16010 7023 7481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_16009 7451 2880 2264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16008 2264 2263 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16007 2264 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16006 7451 2881 2264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_16005 2540 2264 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16004 1999 4161 2398 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16003 2044 2602 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16002 7451 2044 1999 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16001 6283 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_16000 6569 6566 6283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15999 7451 6965 6569 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15998 783 786 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15997 779 787 780 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15996 7451 4161 779 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15995 787 789 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15994 7451 788 789 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15993 7451 785 786 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15992 784 787 783 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15991 782 789 784 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15990 7451 781 782 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15989 781 784 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15988 780 789 781 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15987 7451 780 4161 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15986 4161 780 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15985 7451 1893 1756 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15984 1756 2104 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15983 1756 1896 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15982 7451 6407 1756 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15981 1825 1756 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15980 7451 1852 135 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15979 266 3548 115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15978 115 1852 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15977 115 135 266 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15976 7451 136 115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15975 136 3548 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15974 3391 3389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15973 7451 3997 3390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15972 7451 4577 3392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15971 3419 4577 3391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15970 3390 3392 3419 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15969 3592 3419 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15968 6377 7379 6376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15967 6376 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15966 7451 7335 6377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15965 6375 6377 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15964 4537 4574 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15963 7451 4933 4536 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15962 7451 4577 4578 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15961 4576 4577 4537 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15960 4536 4578 4576 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15959 4572 4576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15958 3613 3870 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15957 7451 3890 3612 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15956 7451 4577 3642 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15955 3641 4577 3613 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15954 3612 3642 3641 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15953 3895 3641 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15952 4219 4217 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15951 7451 4215 4218 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15950 7451 4577 4221 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15949 4220 4577 4219 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15948 4218 4221 4220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15947 4216 4220 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15946 2727 2537 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15945 7451 7162 2727 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15944 5812 5810 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15943 7451 5811 5812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15942 5461 4000 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15941 5461 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15940 7451 6133 5461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15939 7451 6333 5461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15938 4803 4820 4865 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15937 4802 4821 4803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15936 7451 4819 4802 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15935 5815 4865 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15934 2534 2533 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15933 7451 2534 2531 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15932 2532 2866 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15931 7451 2532 2530 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15930 2530 2531 2529 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15929 2529 2534 2528 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15928 2525 3819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_15927 7451 2526 3819 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15926 3819 2526 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15925 2528 2527 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15924 2527 2529 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15923 7451 7500 2527 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15922 2526 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15921 2526 2531 2525 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_15920 2527 2534 2526 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_15919 6983 7508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15918 7451 6983 6987 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15917 6986 6988 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15916 7451 6986 6961 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15915 6961 6987 6985 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15914 6985 6983 6960 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15913 6959 6991 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_15912 7451 6982 6991 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15911 6991 6982 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15910 6960 6984 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15909 6984 6985 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15908 7451 7500 6984 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15907 6982 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15906 6982 6987 6959 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_15905 6984 6983 6982 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_15904 7421 7419 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15903 7422 7470 7421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15902 7451 7420 7422 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15901 5275 4569 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15900 5275 5369 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15899 7451 4568 5275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15898 3734 3817 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15897 7451 3837 3734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15896 7451 3000 1846 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15895 1846 1869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15894 1867 3546 1846 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15893 1845 2095 1867 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15892 1846 1866 1845 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15891 809 3917 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15890 7451 963 808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15889 7451 875 864 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15888 863 875 809 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15887 808 864 863 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15886 968 863 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15885 1156 2435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15884 1155 2853 1156 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15883 7451 2133 1155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15882 5466 7390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15881 5466 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15880 7451 6061 5466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15879 7451 7388 5466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15878 2280 6035 2279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15877 2300 3645 2280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15876 2280 3135 2300 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15875 2279 2926 2280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15874 2279 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15873 7451 5043 2279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15872 516 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15871 778 1085 516 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15870 7451 831 778 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15869 3302 3487 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15868 7451 3409 3302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15867 3300 3302 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15866 2980 5225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15865 3006 4413 2980 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15864 2979 4411 3006 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15863 7451 3005 2979 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15862 3004 3006 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15861 3451 4673 3515 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15860 3514 5000 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15859 7451 3514 3451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15858 1043 2591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15857 7451 3820 1043 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15856 1500 1043 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15855 6428 6954 6469 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15854 6468 6532 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15853 7451 6468 6428 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15852 2555 2926 2556 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15851 2556 3135 2579 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15850 2579 3499 2556 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15849 2555 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15848 7451 5137 2555 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15847 2556 6025 2555 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15846 2576 2579 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15845 1277 1883 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15844 7451 1851 1277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15843 1558 1277 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15842 3945 6846 4006 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15841 4005 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15840 7451 4005 3945 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15839 7451 5718 4073 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15838 4073 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15837 7451 5000 4073 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15836 4149 4073 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15835 1760 2037 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15834 7451 1759 1760 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15833 1973 1760 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15832 2518 2517 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15831 2515 4697 2518 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15830 2516 4695 2515 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15829 7451 2590 2516 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15828 2514 2515 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15827 6826 6828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15826 6821 6829 6822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15825 7451 7481 6821 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15824 6829 6830 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15823 7451 7208 6830 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15822 7451 6825 6828 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15821 6827 6829 6826 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15820 6823 6830 6827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15819 7451 6824 6823 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15818 6824 6827 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15817 6822 6830 6824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15816 7451 6822 7481 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15815 7481 6822 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15814 7087 7086 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15813 7080 7089 7082 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15812 7451 7464 7080 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15811 7089 7088 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15810 7451 7199 7088 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15809 7451 7084 7086 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15808 7085 7089 7087 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15807 7081 7088 7085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15806 7451 7083 7081 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15805 7083 7085 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15804 7082 7088 7083 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15803 7451 7082 7464 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15802 7464 7082 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15801 792 1572 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15800 793 1046 792 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15799 7451 979 793 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15798 6003 6165 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15797 6027 6166 6003 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15796 7451 6125 6027 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15795 7344 7357 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15794 7358 7458 7344 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15793 7451 7420 7358 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15792 5353 5502 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15791 7451 5352 5353 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15790 5500 5411 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15789 7451 7010 5500 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15788 2991 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15787 7451 2591 2991 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15786 761 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15785 760 1465 761 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15784 759 1464 760 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15783 7451 1598 759 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15782 1548 760 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15781 2154 2263 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15780 7451 3023 2154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15779 264 3545 263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15778 263 3549 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15777 7451 3546 264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15776 262 264 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15775 5423 5420 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15774 7451 5421 5423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15773 6446 6631 6423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15772 6423 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15771 7451 7034 6423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15770 6444 6446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15769 6422 7032 6446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15768 6423 7129 6422 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15767 6917 7391 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15766 7451 7384 6917 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15765 5804 7454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15764 5804 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15763 7451 6968 5804 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15762 6021 7379 6001 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15761 6001 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15760 7451 6628 6021 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15759 6160 6021 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15758 5566 5981 5605 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15757 5564 5818 5566 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15756 5565 5819 5564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15755 7451 5815 5565 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_15754 5604 5605 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15753 6530 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15752 6531 6566 6530 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15751 7451 7452 6531 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15750 4568 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15749 4568 4603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15748 7451 4600 4568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15747 7451 6333 4568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15746 7451 6652 6714 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15745 7451 6061 6063 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15744 6714 6063 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15743 2244 2245 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15742 2242 4697 2244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15741 2243 4695 2242 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15740 7451 2442 2243 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15739 2241 2242 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15738 6941 7075 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15737 6940 7255 6941 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15736 7451 7420 6940 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15735 7451 4158 3285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15734 3285 3515 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15733 3356 5043 3285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15732 3284 3922 3356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15731 3285 3925 3284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15730 5252 5690 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15729 5252 5691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15728 7451 5841 5252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15727 2086 2842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15726 2425 2792 2086 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15725 7451 2504 2425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15724 1854 2576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15723 7451 1851 1854 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15722 1852 1854 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15721 7451 6869 6450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15720 6450 6676 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15719 7451 6965 6450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15718 6553 6450 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15717 7451 5093 4510 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15716 4510 4732 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15715 7451 5178 4510 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15714 4585 4510 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15713 7451 5678 5680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15712 5680 5895 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15711 7451 5679 5680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15710 5677 5680 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15709 577 833 543 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15708 543 653 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15707 7451 778 577 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15706 576 577 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15705 1713 2009 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15704 2002 2007 1713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15703 7451 2008 2002 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15702 3258 3738 3257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15701 3257 3665 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15700 7451 3513 3258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15699 3256 3258 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15698 5847 5917 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15697 5848 6058 5847 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15696 7451 5846 5848 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15695 5850 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15694 6010 7379 5850 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15693 7451 7335 6010 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15692 2236 2263 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15691 7451 3023 2236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15690 2292 2236 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15689 7451 7460 7461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15688 7458 7455 7445 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15687 7445 7460 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15686 7445 7461 7458 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15685 7451 7457 7445 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15684 7457 7455 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15683 7254 7387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15682 7289 7513 7254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15681 7451 7287 7289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15680 6390 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15679 6389 6394 6390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15678 7451 6388 6389 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15677 1164 1501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15676 7451 1500 1164 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15675 2543 1164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15674 7451 5989 5990 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15673 5990 5988 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15672 7451 6044 5990 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15671 5987 5990 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15670 6260 6407 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15669 7451 6408 6260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15668 6474 6260 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15667 797 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15666 7451 4376 797 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15665 2880 797 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15664 216 461 199 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15663 199 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15662 7451 511 216 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15661 507 216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15660 7451 1558 1559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15659 1556 1560 1557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15658 1557 1558 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15657 1557 1559 1556 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15656 7451 1555 1557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15655 1555 1560 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15654 7113 7496 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15653 5225 5138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15652 534 533 535 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15651 535 536 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15650 7451 4600 534 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15649 4728 534 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15648 7451 4447 4375 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15647 4375 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15646 4375 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15645 7451 4446 4375 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15644 5994 4375 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15643 3249 3917 3250 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15642 3250 3420 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15641 7451 4823 3249 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15640 3248 3249 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15639 3399 3398 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15638 3393 3401 3394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15637 7451 3696 3393 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15636 3401 3402 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15635 7451 3400 3402 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15634 7451 3695 3398 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15633 3397 3401 3399 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15632 3395 3402 3397 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15631 7451 3396 3395 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15630 3396 3397 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15629 3394 3402 3396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15628 7451 3394 3696 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15627 3696 3394 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15626 7451 7418 7139 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15625 7137 7464 7117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15624 7117 7418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15623 7117 7139 7137 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15622 7451 7135 7117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15621 7135 7464 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15620 4787 5385 5378 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15619 4786 6846 4787 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15618 7451 5467 4786 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15617 2929 4724 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15616 7451 5889 2929 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15615 7201 7379 7202 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15614 7202 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15613 7451 7462 7201 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15612 7261 7201 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15611 3602 3666 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15610 7451 3601 3602 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15609 4172 3602 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15608 2613 2684 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15607 7451 2814 2613 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15606 1428 3545 1429 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15605 1429 1823 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15604 7451 3546 1428 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15603 1427 1428 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15602 7045 7113 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15601 7045 7164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15600 7451 7391 7045 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15599 7451 7114 7045 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15598 5881 5966 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15597 7451 5879 5881 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15596 4034 4574 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15595 7451 6432 4032 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15594 7451 5128 4033 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15593 4035 5128 4034 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15592 4032 4033 4035 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15591 6439 4035 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15590 3607 3870 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15589 7451 6617 3606 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15588 7451 5128 3622 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15587 3623 5128 3607 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15586 3606 3622 3623 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15585 6620 3623 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15584 3277 4217 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15583 7451 3550 3276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15582 7451 5128 3299 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15581 3296 5128 3277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15580 3276 3299 3296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15579 3554 3296 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15578 776 1688 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15577 776 775 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15576 7451 1155 776 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15575 2424 2304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15574 2424 2514 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15573 7451 2383 2424 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15572 5159 5158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15571 7451 5156 5159 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15570 5830 5159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15569 1581 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15568 1581 1707 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15567 7451 4377 1581 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15566 7451 4376 1581 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15565 2678 2679 2677 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15564 2739 5001 2678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15563 2678 5840 2739 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15562 2677 2816 2678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15561 2677 5842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15560 7451 7108 2677 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15559 1624 3742 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15558 1624 1384 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15557 7451 1915 1624 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15556 6774 7049 6724 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15555 6724 6849 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15554 7451 6917 6774 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15553 6773 6774 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15552 7451 7477 7479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15551 7479 7475 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15550 7451 7480 7479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15549 7474 7479 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15548 4771 4979 4358 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15547 4358 5832 4771 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15546 7451 4425 4358 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15545 4789 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15544 4789 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15543 7451 4447 4789 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15542 7451 4446 4789 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15541 7451 4437 4433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15540 4433 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15539 4433 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15538 7451 6333 4433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15537 4995 4433 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15536 7451 2463 2335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15535 2335 2332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15534 7451 2333 2335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15533 3033 2335 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15532 408 479 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15531 406 443 478 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15530 7451 437 406 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15529 443 444 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15528 7451 669 444 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15527 7451 480 479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15526 440 443 408 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15525 407 444 440 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15524 7451 439 407 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15523 439 440 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15522 478 444 439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15521 7451 478 437 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15520 437 478 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15519 7451 765 562 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15518 562 819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15517 7451 1809 562 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15516 696 562 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15515 4688 5275 5351 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15514 4687 4715 4688 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15513 7451 5273 4687 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15512 7451 4158 3920 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15511 7451 4156 3921 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15510 3920 3921 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15509 931 1373 1041 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15508 932 975 931 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15507 7451 1044 932 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15506 7451 4600 1703 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15505 1703 2033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15504 1703 2103 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15503 7451 7162 1703 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15502 2946 1703 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15501 2833 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15500 2860 4669 2833 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15499 7451 2949 2860 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15498 4641 4760 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15497 7451 4762 4641 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15496 4973 5056 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15495 7451 6444 4973 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15494 5576 6538 5626 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15493 5575 5625 5576 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15492 7451 5909 5575 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15491 5703 5720 5846 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15490 5702 6538 5703 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15489 7451 5909 5702 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15488 7451 7486 7374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15487 7377 7488 7347 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15486 7347 7486 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15485 7347 7374 7377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15484 7451 7376 7347 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15483 7376 7488 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15482 7256 7428 7245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15481 7245 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15480 7451 7453 7256 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15479 7255 7256 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15478 5515 4982 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15477 7451 4809 5515 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15476 2878 3178 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15475 7451 3179 2878 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15474 3116 2878 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15473 6851 7387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15472 6851 6912 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15471 7451 7168 6851 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15470 2609 2612 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15469 7451 2608 2609 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15468 5128 2609 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15467 5365 5364 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15466 7451 6099 5365 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15465 7451 1619 1438 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15464 1438 1620 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15463 2220 1834 1438 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15462 1437 3425 2220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15461 1438 1631 1437 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15460 7451 7042 7006 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15459 7006 7109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15458 7044 7384 7006 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15457 7005 7286 7044 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15456 7006 7391 7005 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15455 7451 4215 3942 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15454 3942 4228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15453 5681 3993 3942 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15452 3941 4149 5681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15451 3942 5909 3941 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15450 7381 6907 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15449 7381 6843 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15448 7451 7110 7381 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15447 4928 4927 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15446 7451 4926 4928 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15445 5243 4928 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15444 2695 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15443 2836 2929 2695 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15442 7451 6388 2836 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15441 1362 1837 1322 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15440 1322 2174 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15439 7451 7162 1362 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15438 1431 1362 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15437 2467 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15436 2467 2684 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15435 7451 2880 2467 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15434 7451 2881 2467 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15433 2337 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15432 2337 2263 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15431 7451 2880 2337 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15430 7451 2881 2337 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15429 7451 1021 214 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15428 894 462 198 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15427 198 1021 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15426 198 214 894 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15425 7451 212 198 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15424 212 462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15423 6128 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15422 6128 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15421 7451 5833 6128 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15420 7451 7162 6128 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15419 7451 7418 7259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15418 7259 7464 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15417 7451 7462 7259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15416 7460 7259 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15415 7451 7358 5416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15414 5416 5413 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15413 7451 5804 5416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15412 5505 5416 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15411 2797 4695 2796 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15410 2796 3149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15409 7451 2856 2797 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15408 2795 2797 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15407 2212 2785 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15406 7451 2837 2212 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15405 2287 2212 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15404 271 2696 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15403 7451 1851 271 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15402 272 271 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15401 1972 1971 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15400 7451 2811 1972 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15399 1970 1972 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15398 3098 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15397 3097 4669 3098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15396 7451 3499 3097 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15395 7451 6726 5864 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15394 6014 5860 5849 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15393 5849 6726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15392 5849 5864 6014 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15391 7451 5862 5849 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15390 5862 5860 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15389 7100 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15388 7099 7379 7100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15387 7451 7489 7099 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15386 5404 5448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15385 5402 5447 5443 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15384 7451 5536 5402 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15383 5447 5450 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15382 7451 5449 5450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15381 7451 5535 5448 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15380 5444 5447 5404 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15379 5403 5450 5444 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15378 7451 5442 5403 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15377 5442 5444 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15376 5443 5450 5442 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15375 7451 5443 5536 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15374 5536 5443 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15373 4763 5884 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15372 4762 5885 4763 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15371 7451 5069 4762 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15370 5514 5516 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15369 5509 5517 5510 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15368 7451 7511 5509 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15367 5517 5519 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15366 7451 5518 5519 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15365 7451 5515 5516 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15364 5513 5517 5514 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15363 5512 5519 5513 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15362 7451 5511 5512 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15361 5511 5513 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15360 5510 5519 5511 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15359 7451 5510 7511 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15358 7511 5510 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15357 7451 2300 2089 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15356 2089 2800 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15355 7451 2801 2089 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15354 2088 2089 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15353 2245 2596 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15352 1064 1092 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15351 1284 1091 1064 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15350 7451 1159 1284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15349 3839 4673 3768 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15348 3768 3837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15347 7451 6576 3839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15346 3836 3839 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15345 7014 7078 6994 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15344 6994 7034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15343 7451 7033 6994 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15342 7010 7014 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15341 6993 7032 7014 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15340 6994 7011 6993 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15339 7451 1168 684 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15338 684 1449 5171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15337 4852 4979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15336 2590 3086 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15335 3001 6173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15334 1885 2027 1843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15333 1843 3545 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15332 7451 2029 1885 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15331 3655 1885 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15330 525 528 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15329 521 529 522 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15328 7451 1449 521 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15327 529 530 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15326 7451 598 530 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15325 7451 527 528 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15324 526 529 525 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15323 524 530 526 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15322 7451 523 524 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15321 523 526 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15320 522 530 523 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15319 7451 522 1449 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15318 1449 522 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15317 7451 281 282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15316 282 647 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15315 280 470 282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15314 279 468 280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15313 282 469 279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15312 1817 2661 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15311 1871 2658 1817 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15310 7451 2504 1871 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15309 5817 5746 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15308 1067 2618 1114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15307 1066 1382 1067 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15306 7451 1312 1066 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15305 2125 2149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15304 3142 2154 2125 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15303 7451 2164 3142 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15302 7451 1883 1848 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15301 1848 1880 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15300 2960 1881 1848 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15299 1847 5735 2960 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15298 1848 5734 1847 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15297 7451 6819 6738 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15296 6736 6733 6718 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15295 6718 6819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15294 6718 6738 6736 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15293 7451 6735 6718 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15292 6735 6733 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15291 1595 2542 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15290 1657 1628 1595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15289 1594 2541 1657 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15288 7451 2543 1594 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15287 1627 1657 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15286 5797 5727 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15285 7451 5503 5797 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15284 2385 3389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15283 7451 2664 2384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15282 7451 4106 2387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15281 2386 4106 2385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15280 2384 2387 2386 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15279 2669 2386 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15278 3930 4574 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15277 7451 6804 3929 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15276 7451 4106 3974 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15275 3973 4106 3930 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15274 3929 3974 3973 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15273 6811 3973 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15272 1377 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15271 1377 2591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15270 7451 1976 1377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15269 7451 4376 1377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15268 4539 5385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15267 4595 4594 4539 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15266 4538 6846 4595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15265 7451 4593 4538 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15264 4783 4595 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15263 1834 1833 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15262 7451 7114 1834 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15261 3872 3870 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15260 7451 3868 3869 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15259 7451 4106 3871 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15258 3875 4106 3872 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15257 3869 3871 3875 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15256 3876 3875 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15255 3611 4217 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15254 7451 3774 3610 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15253 7451 4106 3631 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15252 3630 4106 3611 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15251 3610 3631 3630 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15250 3779 3630 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15249 7451 5438 5439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15248 5439 7027 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15247 7451 5604 5439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15246 5670 5439 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15245 5409 5695 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15244 5625 5544 5409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15243 5408 5470 5625 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15242 7451 6714 5408 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15241 7451 7174 7176 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15240 7176 7173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15239 7451 7287 7176 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15238 7243 7176 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15237 6383 6736 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15236 6382 6523 6383 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15235 7451 7420 6382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15234 913 1365 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15233 1363 1501 913 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15232 7451 1500 1363 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15231 2786 3134 2788 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15230 2788 2991 2787 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15229 2787 2995 2788 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15228 2786 2837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15227 7451 2785 2786 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15226 2788 3878 2786 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15225 2784 2787 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15224 7451 771 80 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15223 78 275 79 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15222 79 771 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15221 79 80 78 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15220 7451 77 79 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15219 77 275 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15218 7451 7464 7015 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15217 7015 7418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15216 7015 7454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15215 7451 7462 7015 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15214 7074 7015 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15213 3085 3083 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15212 7451 3084 3085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15211 3636 3085 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15210 7451 1342 1151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15209 1151 1340 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15208 1149 1341 1151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15207 1150 1551 1149 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15206 1151 1741 1150 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15205 3413 3411 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15204 7451 3412 3413 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15203 3410 3413 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15202 5233 5138 4652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15201 4652 5832 5233 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15200 7451 4651 4652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15199 2250 4158 2263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15198 2249 4934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15197 7451 2249 2250 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15196 7451 1974 1975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15195 1975 1973 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15194 7451 2454 1975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15193 4360 1975 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15192 1098 2392 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15191 7451 3820 1098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15190 1366 1098 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15189 1807 2292 1808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15188 1808 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15187 7451 2392 1808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15186 3066 1807 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15185 1806 2287 1807 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15184 1808 2922 1806 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15183 7451 1496 1493 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15182 1493 1825 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15181 1493 2315 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15180 7451 1826 1493 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15179 1565 1493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15178 6418 6461 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15177 6416 6462 6456 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15176 7451 7493 6416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15175 6462 6463 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15174 7451 6693 6463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15173 7451 6466 6461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15172 6458 6462 6418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15171 6417 6463 6458 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15170 7451 6457 6417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15169 6457 6458 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15168 6456 6463 6457 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15167 7451 6456 7493 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15166 7493 6456 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15165 7451 3432 3433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15164 3433 4869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15163 7451 3670 3433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15162 3431 3433 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15161 7451 2431 2426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15160 2426 2429 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15159 2426 2425 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15158 7451 2844 2426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15157 3083 2426 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15156 7451 1149 896 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15155 1075 1809 898 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15154 898 1149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15153 898 896 1075 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15152 7451 897 898 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15151 897 1809 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_15150 5222 5884 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15149 5506 5885 5222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15148 7451 5876 5506 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15147 6278 6304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15146 6276 6303 6296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15145 7451 7475 6276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15144 6303 6305 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15143 7451 6302 6305 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_15142 7451 6594 6304 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15141 6300 6303 6278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15140 6277 6305 6300 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15139 7451 6298 6277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15138 6298 6300 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15137 6296 6305 6298 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_15136 7451 6296 7475 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15135 7475 6296 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15134 4671 7162 4672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15133 4672 4828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15132 7451 6266 4672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15131 4669 4671 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15130 4670 4790 4671 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15129 4672 5016 4670 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15128 4761 4973 4760 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15127 4759 4978 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15126 7451 4759 4761 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15125 4389 4424 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15124 4425 5381 4389 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15123 7451 6386 4425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15122 1091 1041 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15121 7451 1040 1091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15120 7122 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15119 7156 7228 7122 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15118 7451 7481 7156 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15117 1561 1823 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15116 1560 3545 1561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15115 7451 3546 1560 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15114 5092 6408 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15113 5092 5837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15112 7451 6407 5092 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15111 6947 7464 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15110 6947 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15109 7451 6968 6947 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15108 1371 1577 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15107 7451 4158 1371 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15106 1580 1579 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15105 6408 1765 1580 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15104 7451 1906 6408 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15103 7451 2946 1718 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15102 1720 1892 1723 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15101 1719 1753 1720 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15100 1718 2945 1719 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15099 4824 2956 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15098 4824 2988 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15097 7451 2958 4824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15096 1092 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15095 7451 4589 1092 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15094 1764 4597 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15093 7451 1709 1764 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15092 2809 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15091 2861 2946 2809 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15090 7451 5043 2861 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15089 1869 3135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15088 7451 3012 1869 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15087 5392 5467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15086 5720 5466 5392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15085 5391 5544 5720 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15084 7451 5695 5391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_15083 6005 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15082 6037 6394 6005 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15081 7451 6035 6037 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15080 564 563 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15079 564 566 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15078 7451 568 564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15077 7451 2954 2728 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15076 2728 2730 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15075 2728 2743 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15074 7451 2727 2728 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15073 4577 2728 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15072 1989 5882 1988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15071 2023 2949 1989 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15070 1989 3135 2023 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15069 1988 2926 1989 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15068 1988 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15067 7451 5138 1988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15066 7451 5992 5370 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15065 5370 5891 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15064 7451 5889 5370 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15063 5369 5370 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15062 7451 7263 5663 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15061 5663 5662 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15060 7451 6023 5663 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15059 5809 5663 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15058 7451 1075 1078 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15057 1078 1074 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15056 7451 1145 1078 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15055 1267 1078 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15054 7029 7099 7000 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15053 7000 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15052 7451 7034 7000 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15051 7027 7029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15050 6999 7032 7029 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15049 7000 7484 6999 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15048 6398 6400 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15047 7451 6897 6398 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15046 6397 6398 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15045 3634 3633 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15044 7451 3632 3634 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15043 4265 3634 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15042 7451 3240 1649 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15041 1744 1649 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15040 7451 1649 1744 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15039 7451 1649 1744 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15038 1744 1649 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15037 7451 1744 1278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15036 3081 1278 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15035 7451 1278 3081 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15034 7451 1278 3081 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15033 3081 1278 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15032 7451 1744 1745 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15031 3135 1745 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15030 7451 1745 3135 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15029 7451 1745 3135 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15028 3135 1745 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15027 7451 286 287 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15026 390 287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15025 7451 287 390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15024 7451 287 390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15023 390 287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15022 7451 390 189 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15021 2686 189 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15020 7451 189 2686 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15019 7451 189 2686 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15018 2686 189 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15017 7451 390 391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15016 4158 391 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15015 7451 391 4158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15014 7451 391 4158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15013 4158 391 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15012 644 824 645 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15011 645 823 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15010 7451 900 644 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15009 698 644 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_15008 7451 1653 1651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15007 1651 1652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15006 7451 1828 1651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15005 4695 1651 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15004 7451 1376 1048 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15003 1048 1047 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15002 7451 1363 1048 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_15001 1046 1048 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_15000 607 1168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14999 7451 1449 607 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14998 1052 607 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14997 5211 5454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14996 3978 6025 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14995 3770 6804 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14994 4423 4986 4388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14993 4388 5889 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14992 7451 4589 4388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14991 6246 4423 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14990 4387 4987 4423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14989 4388 4984 4387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14988 277 276 278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14987 278 280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14986 7451 512 277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14985 899 277 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14984 4908 5216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14983 4698 5125 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14982 4090 4120 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14981 4088 4123 4115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14980 7451 4113 4088 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14979 4123 4122 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14978 7451 4488 4122 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14977 7451 4119 4120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14976 4118 4123 4090 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14975 4089 4122 4118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14974 7451 4116 4089 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14973 4116 4118 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14972 4115 4122 4116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14971 7451 4115 4113 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14970 4113 4115 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14969 3260 3922 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14968 3259 3925 3260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14967 7451 5216 3259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14966 2108 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14965 2454 2541 2108 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14964 7451 2322 2454 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14963 2182 6333 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14962 2182 1837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14961 7451 4000 2182 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14960 7234 7384 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14959 7234 7356 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14958 7451 7286 7234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14957 5665 6029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14956 5664 6030 5665 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14955 7451 6125 5664 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14954 3281 3326 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14953 7451 4424 3280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14952 7451 4264 3329 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14951 3327 4264 3281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14950 3280 3329 3327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14949 3324 3327 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14948 3762 6894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14947 7451 4718 3761 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14946 7451 4264 3809 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14945 3806 4264 3762 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14944 3761 3809 3806 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14943 3905 3806 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14942 3223 3300 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14941 7451 4991 3222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14940 7451 4264 3225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14939 3224 4264 3223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14938 3222 3225 3224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14937 3568 3224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14936 7451 7098 6838 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14935 6838 6836 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14934 7451 6837 6838 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14933 6892 6838 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14932 7451 7149 6699 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14931 6699 6698 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14930 7451 6696 6699 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14929 6697 6699 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14928 1699 2165 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14927 1699 2241 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14926 7451 2101 1699 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14925 3714 3713 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14924 7451 4431 3711 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14923 7451 4264 3715 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14922 3712 4264 3714 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14921 3711 3715 3712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14920 3953 3712 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14919 1809 4158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14918 1809 2174 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14917 7451 3814 1809 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14916 7451 5690 1809 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14915 4673 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14914 4673 5172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14913 7451 5173 4673 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14912 7451 3742 4673 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14911 7451 6015 5285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14910 5285 5282 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14909 7451 6017 5285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14908 5507 5285 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14907 2663 3156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14906 7451 2662 2663 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14905 3128 2663 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14904 1902 2536 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14903 7451 2602 1902 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14902 2039 1902 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14901 7451 1851 1459 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14900 1459 1876 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14899 1479 1688 1459 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14898 1458 2095 1479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14897 1459 3545 1458 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14896 1861 1860 1842 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14895 1842 2007 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14894 7451 2009 1861 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14893 4984 1861 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14892 7451 7074 7077 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14891 7075 7196 7076 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14890 7076 7074 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14889 7076 7077 7075 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14888 7451 7073 7076 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14887 7073 7196 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14886 1272 1809 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14885 7451 1271 1272 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14884 1270 1272 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14883 3172 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14882 7451 6980 3172 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14881 3170 3172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14880 2857 3232 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14879 7451 2948 2857 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14878 2856 2857 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14877 7451 777 711 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14876 711 778 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14875 7451 776 711 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14874 709 711 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14873 416 468 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14872 515 469 416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14871 7451 470 515 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14870 7451 4603 1774 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14869 1774 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14868 7451 6133 1774 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14867 1771 1774 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14866 2271 2313 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14865 2269 2312 2307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14864 7451 2596 2269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14863 2312 2314 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14862 7451 2672 2314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14861 7451 2597 2313 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14860 2309 2312 2271 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14859 2270 2314 2309 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14858 7451 2308 2270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14857 2308 2309 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14856 2307 2314 2308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14855 7451 2307 2596 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14854 2596 2307 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14853 7451 1384 1241 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14852 1241 1915 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14851 7451 3742 1241 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14850 1211 1241 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14849 6831 7466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14848 6831 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14847 7451 6968 6831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14846 7451 5378 3445 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14845 3446 5541 3729 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14844 3444 3456 3446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14843 3445 5377 3444 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14842 4505 4504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14841 4651 5381 4505 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14840 7451 6386 4651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14839 1765 4597 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14838 7451 1624 1765 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14837 7451 7390 6853 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14836 6853 7388 6854 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14835 6852 6854 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14834 6393 6576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14833 6393 6336 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14832 7451 6112 6393 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14831 5571 5617 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14830 6315 5616 5571 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14829 7451 5889 6315 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14828 1456 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_14827 1810 1465 1456 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_14826 1455 1598 1810 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_14825 7451 1464 1455 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_14824 1881 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14823 1881 1723 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14822 7451 1430 1881 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14821 6550 7074 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14820 7451 7453 6550 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14819 6518 6550 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14818 4366 6600 4912 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14817 4365 4364 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14816 7451 4365 4366 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14815 7451 4296 2821 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14814 2821 6339 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14813 7451 2820 2821 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14812 2819 2821 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14811 7451 7242 6203 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14810 6203 6202 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14809 7451 7111 6203 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14808 6272 6203 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14807 2011 2007 1984 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14806 1984 2009 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14805 7451 2008 2011 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14804 2081 2011 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14803 7451 6382 5968 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14802 5968 5967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14801 7451 6102 5968 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14800 5966 5968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14799 3617 3958 3639 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14798 3618 6030 3617 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14797 7451 3957 3618 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14796 4211 3639 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14795 5947 5949 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14794 5943 5950 5944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14793 7451 7453 5943 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14792 5950 5951 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14791 7451 6231 5951 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14790 7451 5954 5949 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14789 5948 5950 5947 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14788 5946 5951 5948 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14787 7451 5945 5946 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14786 5945 5948 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14785 5944 5951 5945 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14784 7451 5944 7453 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14783 7453 5944 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14782 646 2371 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14781 7451 1851 646 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14780 771 646 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14779 6647 6644 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14778 7451 6840 6647 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14777 6646 6647 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14776 1831 2041 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14775 7451 1830 1831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14774 1832 1831 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14773 1829 2102 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14772 7451 4773 1829 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14771 1828 1829 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14770 7451 6902 6904 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14769 6904 7320 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14768 7451 7039 6904 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14767 6901 6904 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14766 5561 5596 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14765 5559 5595 5589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14764 7451 6676 5559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14763 5595 5597 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14762 7451 5594 5597 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14761 7451 5881 5596 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14760 5591 5595 5561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14759 5560 5597 5591 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14758 7451 5590 5560 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14757 5590 5591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14756 5589 5597 5590 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14755 7451 5589 6676 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14754 6676 5589 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14753 2808 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14752 3009 2946 2808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14751 7451 5274 3009 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14750 5049 5052 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14749 5044 5053 5046 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14748 7451 5045 5044 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14747 5053 5054 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14746 7451 5270 5054 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14745 7451 5051 5052 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14744 5050 5053 5049 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14743 5048 5054 5050 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14742 7451 5047 5048 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14741 5047 5050 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14740 5046 5054 5047 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14739 7451 5046 5045 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14738 5045 5046 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14737 7451 1825 1827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14736 1827 2315 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14735 7451 1826 1827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14734 2288 1827 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14733 1242 1908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14732 7451 1915 1242 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14731 1579 1242 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14730 4197 6388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14729 5555 5554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14728 7451 5555 5553 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14727 5552 5848 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14726 7451 5552 5551 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14725 5551 5553 5550 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14724 5550 5555 5549 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14723 5546 6061 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14722 7451 5547 6061 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14721 6061 5547 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14720 5549 5548 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14719 5548 5550 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14718 7451 7500 5548 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14717 5547 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14716 5547 5553 5546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14715 5548 5555 5547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14714 5606 5523 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14713 3705 5887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14712 5981 6187 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14711 6006 6111 6041 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14710 6040 6039 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14709 7451 6040 6006 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14708 2116 2120 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14707 2112 2119 2113 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14706 7451 2111 2112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14705 2119 2121 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14704 7451 2553 2121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14703 7451 2118 2120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14702 2117 2119 2116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14701 2115 2121 2117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14700 7451 2114 2115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14699 2114 2117 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14698 2113 2121 2114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14697 7451 2113 2111 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14696 2111 2113 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14695 3620 3663 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14694 3830 6340 3620 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14693 7451 3737 3830 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14692 7451 4934 672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14691 672 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14690 672 1449 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14689 7451 4376 672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14688 1908 672 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14687 4255 6392 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14686 4379 6894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14685 5051 4401 4379 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14684 7451 4629 5051 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14683 5226 7164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14682 7451 7286 5226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14681 7211 7210 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14680 7212 7270 7211 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14679 7451 7420 7212 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14678 6319 6318 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14677 7451 6386 6319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14676 6836 6319 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14675 1987 2088 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14674 3957 2153 1987 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14673 7451 2018 3957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14672 6534 6912 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14671 7451 7168 6534 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14670 5084 5083 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14669 7451 5082 5084 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14668 5678 5084 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14667 7252 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14666 7433 7383 7252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14665 7451 7453 7433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14664 7451 4427 4225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14663 4225 4231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14662 4225 4370 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14661 7451 4224 4225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14660 4364 4225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14659 7253 7388 7286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14658 7285 7390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14657 7451 7285 7253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14656 1967 2101 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14655 1967 2023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14654 7451 2241 1967 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14653 7451 2165 1967 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14652 7451 3660 3662 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14651 3662 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14650 7451 4724 3662 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14649 3659 3662 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14648 513 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14647 512 1187 513 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14646 7451 906 512 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14645 3076 3074 3075 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14644 3072 3069 3076 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14643 3073 3070 3072 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14642 7451 3071 3073 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14641 6169 3075 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14640 2388 2743 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14639 7451 6344 2388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14638 2676 2388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14637 2654 2652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14636 7451 2653 2654 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14635 2655 2654 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14634 2372 2926 2374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14633 2374 3081 2373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14632 2373 3226 2374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14631 2372 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14630 7451 5274 2372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14629 2374 5887 2372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14628 2371 2373 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14627 1962 2842 1961 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14626 1961 2792 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14625 7451 2371 1962 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14624 2149 1962 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14623 7451 6914 6396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14622 6396 6529 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14621 6698 6392 6396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14620 6395 6393 6698 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14619 6396 6394 6395 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14618 7451 2591 1101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14617 1101 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14616 7451 2881 1101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14615 1368 1101 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14614 7451 1771 1596 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14613 1596 1838 1632 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14612 4351 4353 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14611 4348 4354 4347 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14610 7451 5882 4348 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14609 4354 4355 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14608 7451 4488 4355 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14607 7451 4416 4353 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14606 4352 4354 4351 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14605 4349 4355 4352 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14604 7451 4350 4349 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14603 4350 4352 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14602 4347 4355 4350 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14601 7451 4347 5882 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14600 5882 4347 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14599 7451 1700 958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14598 958 1968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14597 958 1435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14596 7451 4368 958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14595 960 958 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14594 7451 1700 1038 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14593 1038 1968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14592 1038 1435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14591 7451 1688 1038 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14590 1037 1038 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14589 1578 1709 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14588 1577 1624 1578 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14587 7451 4597 1577 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14586 7451 4448 4004 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14585 4004 4441 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14584 4004 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14583 7451 4934 4004 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14582 5691 4004 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14581 5158 5055 4775 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14580 4775 5832 5158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14579 7451 4862 4775 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14578 6964 7428 6943 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14577 6943 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14576 7451 6965 6964 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14575 6942 6964 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14574 6882 7475 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14573 6882 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14572 7451 6968 6882 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14571 6151 6519 6137 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14570 6137 7034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14569 7451 7033 6137 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14568 6150 6151 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14567 6136 7032 6151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14566 6137 6291 6136 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14565 7451 576 224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14564 907 225 201 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14563 201 576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14562 201 224 907 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14561 7451 222 201 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14560 222 225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14559 2290 3135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14558 7451 3499 2290 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14557 7242 4937 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14556 7242 4938 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14555 7451 6135 7242 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14554 6252 6648 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14553 7451 6839 6252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14552 6386 6252 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14551 6897 7481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14550 6897 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14549 7451 6980 6897 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14548 2281 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14547 2304 2929 2281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14546 7451 6173 2304 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14545 1563 2292 1564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14544 1564 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14543 7451 2392 1564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14542 1965 1563 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14541 1562 2159 1563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14540 1564 2095 1562 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14539 2750 6339 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14538 7451 2820 2750 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14537 2751 2750 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14536 7451 2708 648 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14535 648 1037 649 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14534 647 649 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14533 930 4934 2591 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14532 974 2686 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14531 7451 974 930 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14530 3517 5623 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14529 7451 6333 3517 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14528 3516 3517 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14527 6520 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14526 6519 7379 6520 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14525 7451 7452 6519 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14524 7451 3957 3936 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14523 3936 3958 3983 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14522 6029 3983 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14521 7451 4437 1325 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14520 1325 1368 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14519 1369 1365 1325 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14518 1324 1366 1369 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14517 1325 1500 1324 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14516 3242 5378 3243 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14515 3241 5377 3242 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14514 7451 5541 3241 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_14513 3240 3243 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14512 7451 126 25 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14511 370 78 8 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14510 8 126 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14509 8 25 370 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14508 7451 23 8 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14507 23 78 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14506 7451 3347 3344 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14505 3344 4372 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14504 3344 3348 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14503 7451 3343 3344 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14502 3346 3344 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14501 3318 3571 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14500 7451 3318 3319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14499 3317 3315 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14498 7451 3317 3272 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14497 3272 3319 3314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14496 3314 3318 3271 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14495 3270 4502 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14494 7451 3311 4502 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14493 4502 3311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14492 3271 3312 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14491 3312 3314 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14490 7451 5100 3312 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14489 3311 5100 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14488 3311 3319 3270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14487 3312 3318 3311 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14486 7451 5994 3923 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14485 3923 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14484 7451 5000 3923 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14483 3922 3923 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14482 510 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14481 902 2134 510 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14480 7451 509 902 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14479 7451 790 791 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14478 791 2816 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14477 7451 3023 791 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14476 975 791 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14475 7451 1954 1639 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14474 1639 1810 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14473 7451 1809 1639 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14472 1860 1639 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14471 1460 2424 1461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14470 1461 1699 1483 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14469 1483 2504 1461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14468 1460 2789 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14467 7451 2416 1460 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14466 1461 2502 1460 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14465 2090 1483 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14464 7451 7381 7382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14463 7490 7382 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14462 7451 7382 7490 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14461 7451 7382 7490 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14460 7490 7382 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14459 7451 7490 7281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14458 7280 7281 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14457 7451 7281 7280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14456 7451 7281 7280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14455 7280 7281 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14454 7451 7490 7492 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14453 7491 7492 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14452 7451 7492 7491 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14451 7451 7492 7491 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14450 7491 7492 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14449 7084 6876 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14448 7451 6681 7084 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14447 7451 1037 806 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14446 806 2300 831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14445 7451 3820 671 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14444 671 3352 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14443 7451 4376 671 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14442 1049 671 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14441 3913 3997 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14440 3710 4113 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14439 4916 5043 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14438 5543 7390 5542 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14437 5542 7388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14436 7451 7384 5543 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14435 5541 5543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14434 7451 2810 2382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14433 2382 2381 2383 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14432 7451 5842 5843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14431 5843 7108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14430 5902 5840 5843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14429 5839 5841 5902 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14428 5843 6133 5839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14427 7451 1264 311 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14426 310 311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14425 7451 311 310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14424 7451 311 310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14423 310 311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14422 7451 1264 359 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14421 358 359 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14420 7451 359 358 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14419 7451 359 358 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14418 358 359 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14417 7451 1264 361 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14416 360 361 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14415 7451 361 360 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14414 7451 361 360 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14413 360 361 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14412 7451 1264 317 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14411 316 317 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14410 7451 317 316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14409 7451 317 316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14408 316 317 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14407 7451 1264 367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14406 366 367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14405 7451 367 366 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14404 7451 367 366 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14403 366 367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14402 7451 1264 369 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14401 368 369 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14400 7451 369 368 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14399 7451 369 368 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14398 368 369 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14397 7451 1264 1219 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14396 1180 1219 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14395 7451 1219 1180 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14394 7451 1219 1180 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14393 1180 1219 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14392 7424 7466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14391 6629 6628 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14390 5574 5912 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14389 6195 5623 5574 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14388 7451 6333 6195 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14387 6582 6599 7032 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14386 6581 6848 6582 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14385 7451 6600 6581 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14384 2791 2842 2790 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14383 2790 2792 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14382 7451 2789 2791 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14381 3069 2791 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14380 7168 7236 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14379 7451 7287 7168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14378 7451 1264 1254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14377 1253 1254 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14376 7451 1254 1253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14375 7451 1254 1253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14374 1253 1254 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14373 7451 1264 1256 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14372 1255 1256 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14371 7451 1256 1255 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14370 7451 1256 1255 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14369 1255 1256 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14368 7451 1264 1222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14367 1185 1222 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14366 7451 1222 1185 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14365 7451 1222 1185 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14364 1185 1222 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14363 7451 1264 1262 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14362 1261 1262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14361 7451 1262 1261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14360 7451 1262 1261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14359 1261 1262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14358 7451 1264 1265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14357 1263 1265 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14356 7451 1265 1263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14355 7451 1265 1263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14354 1263 1265 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14353 7451 1281 321 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14352 320 321 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14351 7451 321 320 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14350 7451 321 320 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14349 320 321 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14348 7451 1281 375 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14347 374 375 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14346 7451 375 374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14345 7451 375 374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14344 374 375 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14343 7451 1281 377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14342 376 377 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14341 7451 377 376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14340 7451 377 376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14339 376 377 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14338 5015 5554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14337 7451 5015 5013 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14336 5014 5012 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14335 7451 5014 4958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14334 4958 5013 5010 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14333 5010 5015 4957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14332 4956 7235 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14331 7451 5006 7235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14330 7235 5006 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14329 4957 5008 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14328 5008 5010 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14327 7451 7500 5008 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14326 5006 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14325 5006 5013 4956 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14324 5008 5015 5006 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_14323 511 827 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14322 7451 564 511 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14321 1830 7114 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14320 1830 1837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14319 7451 4158 1830 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14318 1095 1363 1060 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14317 1060 2255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14316 7451 1449 1095 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14315 1203 1095 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14314 3670 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14313 7451 5001 3670 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14312 5695 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14311 7451 6061 5695 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14310 6820 6869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14309 7451 6965 6820 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14308 6819 6820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14307 6340 3159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14306 6340 3303 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14305 7451 3160 6340 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14304 7451 3326 6340 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14303 6273 6272 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14302 7451 6271 6273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14301 6341 6273 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14300 7361 7418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14299 7451 7464 7361 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14298 7413 7361 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14297 7451 1281 327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14296 326 327 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14295 7451 327 326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14294 7451 327 326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14293 326 327 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14292 7451 1281 383 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14291 382 383 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14290 7451 383 382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14289 7451 383 382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14288 382 383 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14287 7451 1281 385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14286 384 385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14285 7451 385 384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14284 7451 385 384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14283 384 385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14282 7451 1281 1224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14281 1190 1224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14280 7451 1224 1190 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14279 7451 1224 1190 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14278 1190 1224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14277 7451 1281 1274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14276 1273 1274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14275 7451 1274 1273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14274 7451 1274 1273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14273 1273 1274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14272 7451 1281 1276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14271 1275 1276 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14270 7451 1276 1275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14269 7451 1276 1275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14268 1275 1276 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14267 7451 1281 1227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14266 1196 1227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14265 7451 1227 1196 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14264 7451 1227 1196 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14263 1196 1227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14262 7451 5752 5733 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14261 6739 5733 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14260 7451 5733 6739 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14259 7451 5733 6739 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14258 6739 5733 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14257 7451 5752 5753 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14256 6771 5753 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14255 7451 5753 6771 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14254 7451 5753 6771 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14253 6771 5753 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14252 7451 3717 3718 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14251 5752 3718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14250 7451 3718 5752 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14249 7451 3718 5752 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14248 5752 3718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14247 3470 1341 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14246 3470 1020 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14245 7451 1025 3470 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14244 1257 1341 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14243 1257 1216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14242 7451 1634 1257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14241 2617 2819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14240 7451 3248 2617 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14239 2884 2617 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14238 7451 5830 5831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14237 5831 7031 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14236 7451 5828 5831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14235 5829 5831 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14234 7451 1412 736 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14233 735 736 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14232 7451 736 735 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14231 7451 736 735 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14230 735 736 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14229 7451 735 673 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14228 5100 673 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14227 7451 673 5100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14226 7451 673 5100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14225 5100 673 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14224 7451 735 299 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14223 7500 299 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14222 7451 299 7500 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14221 7451 299 7500 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14220 7500 299 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14219 1986 2658 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14218 2016 2661 1986 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14217 7451 2133 2016 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14216 7451 4568 4281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14215 4281 4569 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14214 7451 4773 4281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14213 4427 4281 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14212 7451 1281 1280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14211 1279 1280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14210 7451 1280 1279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14209 7451 1280 1279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14208 1279 1280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14207 7451 1281 1283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14206 1282 1283 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14205 7451 1283 1282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14204 7451 1283 1282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14203 1282 1283 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14202 7451 3210 2138 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14201 2137 2138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14200 7451 2138 2137 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14199 7451 2138 2137 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14198 2137 2138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14197 7451 3210 2214 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14196 2213 2214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14195 7451 2214 2213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14194 7451 2214 2213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14193 2213 2214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14192 7451 3210 2216 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14191 2215 2216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14190 7451 2216 2215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14189 7451 2216 2215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14188 2215 2216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14187 7451 3210 2146 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14186 2145 2146 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14185 7451 2146 2145 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14184 7451 2146 2145 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14183 2145 2146 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14182 7451 3210 2225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14181 2224 2225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14180 7451 2225 2224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14179 7451 2225 2224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14178 2224 2225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14177 7451 3210 2227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14176 2226 2227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14175 7451 2227 2226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14174 7451 2227 2226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14173 2226 2227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14172 7451 7466 7367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14171 7367 7477 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14170 7367 7475 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14169 7451 7480 7367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14168 7418 7367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14167 1030 1029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14166 7451 1145 1030 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14165 1034 1030 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14164 2961 3663 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14163 3338 2960 2961 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14162 7451 3256 3338 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14161 7451 7164 5219 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14160 5219 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14159 5218 5216 5219 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14158 5217 5275 5218 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14157 5219 5273 5217 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14156 2439 2862 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14155 7451 2589 2439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14154 2801 2439 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14153 4078 4157 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14152 7451 4377 4078 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14151 4077 4078 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14150 7451 3472 3474 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14149 3474 3469 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14148 7451 3470 3474 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14147 6894 3474 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14146 3557 3559 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14145 3551 3560 3552 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14144 7451 3550 3551 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14143 3560 3561 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14142 7451 3558 3561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14141 7451 3554 3559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14140 3556 3560 3557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14139 3555 3561 3556 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14138 7451 3553 3555 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14137 3553 3556 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14136 3552 3561 3553 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14135 7451 3552 3550 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14134 3550 3552 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14133 976 1384 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14132 7451 2881 976 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14131 1365 976 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14130 769 903 770 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14129 770 768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14128 7451 1732 769 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14127 767 769 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14126 7451 7432 7434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14125 7434 7433 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14124 7451 7430 7434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14123 7431 7434 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14122 1995 2039 2041 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14121 1994 2040 1995 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14120 7451 2456 1994 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14119 7451 2880 2680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14118 2680 2684 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14117 2680 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14116 7451 2881 2680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14115 2679 2680 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14114 6415 6440 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14113 6413 6441 6434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14112 7451 6432 6413 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14111 6441 6442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14110 7451 6622 6442 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_14109 7451 6439 6440 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14108 6436 6441 6415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14107 6414 6442 6436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14106 7451 6435 6414 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14105 6435 6436 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14104 6434 6442 6435 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_14103 7451 6434 6432 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14102 6432 6434 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14101 6013 6010 5999 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14100 5999 7034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14099 7451 7033 5999 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14098 6009 6013 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14097 5998 7032 6013 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14096 5999 6226 5998 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14095 5741 5670 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14094 7451 5671 5741 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14093 2738 2540 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14092 7451 2684 2738 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14091 1812 6175 1811 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14090 2141 3646 1812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14089 1812 3081 2141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14088 1811 2926 1812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14087 1811 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14086 7451 4834 1811 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14085 7451 1733 1472 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14084 2082 1468 1457 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14083 1457 1733 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14082 1457 1472 2082 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14081 7451 1469 1457 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14080 1469 1468 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_14079 7451 3264 3188 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14078 3187 3188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14077 7451 3188 3187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14076 7451 3188 3187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14075 3187 3188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14074 7451 3264 3262 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14073 3261 3262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14072 7451 3262 3261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14071 7451 3262 3261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14070 3261 3262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14069 7451 3264 3265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14068 3263 3265 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14067 7451 3265 3263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14066 7451 3265 3263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14065 3263 3265 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14064 7451 2746 865 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14063 1295 865 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14062 7451 865 1295 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14061 7451 865 1295 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14060 1295 865 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14059 193 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14058 193 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14057 7451 3346 193 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14056 2889 7108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14055 2889 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14054 7451 3346 2889 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14053 6874 7428 6855 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14052 6855 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14051 7451 7454 6874 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14050 7357 6874 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14049 6741 7481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14048 6741 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14047 7451 6968 6741 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14046 2133 1430 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14045 7451 1466 2133 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14044 643 699 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14043 765 698 643 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14042 7451 1341 765 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14041 1740 3135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14040 7451 2949 1740 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14039 2097 2946 2098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14038 2098 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14037 7451 4979 2097 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14036 2381 2097 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_14035 162 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14034 162 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14033 7451 3346 162 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14032 338 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14031 338 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14030 7451 3346 338 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14029 7451 2746 874 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14028 1310 874 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14027 7451 874 1310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14026 7451 874 1310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14025 1310 874 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14024 7451 2746 2726 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14023 3246 2726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14022 7451 2726 3246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14021 7451 2726 3246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14020 3246 2726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14019 7451 2746 2747 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14018 3264 2747 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14017 7451 2747 3264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14016 7451 2747 3264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14015 3264 2747 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14014 1111 2880 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14013 1111 1051 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14012 7451 4442 1111 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14011 875 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14010 875 1292 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14009 7451 4600 875 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14008 2406 2435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14007 2431 2853 2406 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14006 7451 2789 2431 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14005 6336 6333 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14004 6336 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14003 7451 7108 6336 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_14002 5395 6168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14001 5655 6169 5395 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_14000 7451 5876 5655 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13999 7451 5280 4194 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13998 4193 4194 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13997 7451 4194 4193 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13996 7451 4194 4193 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13995 4193 4194 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13994 7451 5280 4246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13993 4245 4246 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13992 7451 4246 4245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13991 7451 4246 4245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13990 4245 4246 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13989 7451 5280 4248 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13988 4247 4248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13987 7451 4248 4247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13986 7451 4248 4247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13985 4247 4248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13984 7451 5280 4199 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13983 4198 4199 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13982 7451 4199 4198 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13981 7451 4199 4198 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13980 4198 4199 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13979 7451 5280 4252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13978 4251 4252 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13977 7451 4252 4251 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13976 7451 4252 4251 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13975 4251 4252 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13974 7451 5280 4253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13973 4638 4253 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13972 7451 4253 4638 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13971 7451 4253 4638 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13970 4638 4253 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13969 7451 5280 5213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13968 5212 5213 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13967 7451 5213 5212 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13966 7451 5213 5212 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13965 5212 5213 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13964 7451 5243 5244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13963 5244 6888 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13962 7451 5241 5244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13961 5242 5244 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13960 6840 7489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13959 6840 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13958 7451 6980 6840 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13957 2436 2853 2407 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13956 2407 2435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13955 7451 2433 2436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13954 2434 2436 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13953 4801 4861 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13952 4862 5381 4801 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13951 7451 6839 4862 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13950 3161 3160 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13949 7451 3159 3161 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13948 3387 3161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13947 7451 190 192 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13946 191 192 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13945 7451 192 191 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13944 7451 192 191 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13943 191 192 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13942 7451 191 31 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13941 7042 31 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13940 7451 31 7042 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13939 7451 31 7042 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13938 7042 31 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13937 7451 191 159 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13936 5841 159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13935 7451 159 5841 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13934 7451 159 5841 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13933 5841 159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13932 7451 5280 5269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13931 5268 5269 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13930 7451 5269 5268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13929 7451 5269 5268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13928 5268 5269 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13927 7451 5280 5271 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13926 5270 5271 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13925 7451 5271 5270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13924 7451 5271 5270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13923 5270 5271 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13922 7451 5280 5221 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13921 5220 5221 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13920 7451 5221 5220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13919 7451 5221 5220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13918 5220 5221 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13917 7451 5280 5279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13916 5278 5279 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13915 7451 5279 5278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13914 7451 5279 5278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13913 5278 5279 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13912 7451 5280 5281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13911 5584 5281 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13910 7451 5281 5584 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13909 7451 5281 5584 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13908 5584 5281 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13907 7451 5296 4205 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13906 4204 4205 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13905 7451 4205 4204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13904 7451 4205 4204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13903 4204 4205 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13902 7451 5296 4259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13901 4258 4259 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13900 7451 4259 4258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13899 7451 4259 4258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13898 4258 4259 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13897 7451 5296 4260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13896 4488 4260 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13895 7451 4260 4488 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13894 7451 4260 4488 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13893 4488 4260 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13892 3800 4561 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13891 7451 3800 3799 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13890 3798 3797 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13889 7451 3798 3751 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13888 3751 3799 3795 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13887 3795 3800 3750 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13886 3749 4861 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13885 7451 3791 4861 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13884 4861 3791 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13883 3750 3792 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13882 3792 3795 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13881 7451 7500 3792 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13880 3791 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13879 3791 3799 3749 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13878 3792 3800 3791 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13877 6287 6344 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13876 6614 6410 6287 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13875 7451 6491 6614 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13874 4521 5385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13873 4519 4602 4521 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13872 4520 4518 4519 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13871 7451 4593 4520 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13870 4517 4519 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13869 7451 2754 1982 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13868 1981 1982 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13867 7451 1982 1981 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13866 7451 1982 1981 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13865 1981 1982 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13864 7451 1981 1388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13863 5690 1388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13862 7451 1388 5690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13861 7451 1388 5690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13860 5690 1388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13859 7451 1981 1710 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13858 7162 1710 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13857 7451 1710 7162 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13856 7451 1710 7162 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13855 7162 1710 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13854 7451 1981 1582 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13853 6333 1582 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13852 7451 1582 6333 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13851 7451 1582 6333 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13850 6333 1582 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13849 7451 1981 1451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13848 7114 1451 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13847 7451 1451 7114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13846 7451 1451 7114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13845 7114 1451 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13844 5962 5961 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13843 5956 5964 5955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13842 7451 7462 5956 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13841 5964 5963 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13840 7451 6302 5963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13839 7451 5960 5961 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13838 5958 5964 5962 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13837 5959 5963 5958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13836 7451 5957 5959 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13835 5957 5958 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13834 5955 5963 5957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13833 7451 5955 7462 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13832 7462 5955 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13831 3723 4360 3725 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13830 3725 3724 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13829 7451 6397 3723 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13828 3722 3723 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13827 2321 2319 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13826 7451 2958 2321 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13825 2318 2321 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13824 2832 3710 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13823 2853 4695 2832 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13822 7451 3145 2853 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13821 1450 4158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13820 7451 1449 1450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13819 1707 1450 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13818 7451 5296 4214 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13817 4213 4214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13816 7451 4214 4213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13815 7451 4214 4213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13814 4213 4214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13813 7451 5296 4269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13812 4268 4269 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13811 7451 4269 4268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13810 7451 4269 4268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13809 4268 4269 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13808 7451 5296 4270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13807 4561 4270 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13806 7451 4270 4561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13805 7451 4270 4561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13804 4561 4270 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13803 7451 5296 5224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13802 5223 5224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13801 7451 5224 5223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13800 7451 5224 5223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13799 5223 5224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13798 7451 5296 5289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13797 5288 5289 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13796 7451 5289 5288 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13795 7451 5289 5288 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13794 5288 5289 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13793 7451 5296 5290 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13792 5594 5290 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13791 7451 5290 5594 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13790 7451 5290 5594 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13789 5594 5290 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13788 7451 5296 5231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13787 5232 5231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13786 7451 5231 5232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13785 7451 5231 5232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13784 5232 5231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13783 5558 5586 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13782 5556 5585 5578 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13781 7451 7335 5556 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13780 5585 5587 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13779 7451 5584 5587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13778 7451 5581 5586 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13777 5582 5585 5558 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13776 5557 5587 5582 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13775 7451 5579 5557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13774 5579 5582 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13773 5578 5587 5579 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13772 7451 5578 7335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13771 7335 5578 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13770 484 4728 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13769 7451 6266 484 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13768 494 484 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13767 3286 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13766 3432 7108 3286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13765 7451 6332 3432 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13764 4902 4905 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13763 4898 4904 4899 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13762 7451 5350 4898 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13761 4904 4906 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13760 7451 5584 4906 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13759 7451 5353 4905 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13758 4903 4904 4902 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13757 4901 4906 4903 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13756 7451 4900 4901 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13755 4900 4903 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13754 4899 4906 4900 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13753 7451 4899 5350 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13752 5350 4899 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13751 7473 7475 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13750 1587 2926 1588 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13749 1588 3135 1646 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13748 1646 2949 1588 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13747 1587 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13746 7451 5138 1587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13745 1588 5882 1587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13744 1883 1646 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13743 7451 5296 5295 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13742 5294 5295 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13741 7451 5295 5294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13740 7451 5295 5294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13739 5294 5295 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13738 7451 5296 5297 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13737 5518 5297 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13736 7451 5297 5518 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13735 7451 5297 5518 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13734 5518 5297 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13733 7451 7194 6149 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13732 6148 6149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13731 7451 6149 6148 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13730 7451 6149 6148 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13729 6148 6149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13728 7451 7194 6223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13727 6222 6223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13726 7451 6223 6222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13725 7451 6223 6222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13724 6222 6223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13723 7451 7194 6224 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13722 6622 6224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13721 7451 6224 6622 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13720 7451 6224 6622 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13719 6622 6224 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13718 7451 7194 6155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13717 6154 6155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13716 7451 6155 6154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13715 7451 6155 6154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13714 6154 6155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13713 7451 7194 6230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13712 6229 6230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13711 7451 6230 6229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13710 7451 6230 6229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13709 6229 6230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13708 7451 7194 6232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13707 6231 6232 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13706 7451 6232 6231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13705 7451 6232 6231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13704 6231 6232 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13703 7513 7512 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13702 5860 7335 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13701 4282 4782 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13700 4919 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13699 5075 5273 4919 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13698 7451 6388 5075 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13697 3207 3214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13696 3484 3212 3207 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13695 7451 3475 3484 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13694 2286 2841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13693 7451 2836 2286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13692 7094 7481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13691 1631 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13690 7451 1976 1631 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13689 3667 3119 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13688 7451 3266 3667 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13687 5376 5992 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13686 7451 5891 5376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13685 6294 7379 6275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13684 6275 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13683 7451 7452 6294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13682 6293 6294 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13681 7316 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13680 7451 7493 7331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13679 7330 7494 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13678 7451 7330 7316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13677 7316 7331 7329 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13676 7329 7494 7316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13675 7315 7329 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13674 7451 7329 7315 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13673 7451 7194 7125 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13672 7124 7125 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13671 7451 7125 7124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13670 7451 7125 7124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13669 7124 7125 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13668 7451 7194 7188 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13667 7187 7188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13666 7451 7188 7187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13665 7451 7188 7187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13664 7187 7188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13663 7451 7194 7190 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13662 7189 7190 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13661 7451 7190 7189 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13660 7451 7190 7189 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13659 7189 7190 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13658 7451 7194 7127 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13657 7126 7127 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13656 7451 7127 7126 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13655 7451 7127 7126 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13654 7126 7127 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13653 7451 7194 7192 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13652 7191 7192 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13651 7451 7192 7191 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13650 7451 7192 7191 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13649 7191 7192 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13648 7451 7194 7195 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13647 7193 7195 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13646 7451 7195 7193 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13645 7451 7195 7193 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13644 7193 7195 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13643 7451 7207 6164 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13642 6163 6164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13641 7451 6164 6163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13640 7451 6164 6163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13639 6163 6164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13638 7509 7508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13637 7451 7509 7510 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13636 7507 7505 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13635 7451 7507 7450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13634 7450 7510 7504 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13633 7504 7509 7449 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13632 7448 7496 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13631 7451 7499 7496 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13630 7496 7499 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13629 7449 7502 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13628 7502 7504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13627 7451 7500 7502 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13626 7499 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13625 7499 7510 7448 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13624 7502 7509 7499 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13623 6427 6600 6467 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13622 6426 6599 6427 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13621 7451 6848 6426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13620 7420 6467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13619 2969 3263 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13618 7451 2969 2970 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13617 2967 2973 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13616 7451 2967 2968 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13615 2968 2970 2965 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13614 2965 2969 2966 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13613 2962 3814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13612 7451 2963 3814 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13611 3814 2963 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13610 2966 2964 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13609 2964 2965 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13608 7451 7500 2964 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13607 2963 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13606 2963 2970 2962 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13605 2964 2969 2963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13604 906 2371 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13603 7451 1851 906 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13602 7451 4376 340 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13601 7451 4161 194 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13600 340 194 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13599 6267 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13598 7451 6266 6267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13597 7451 7207 6238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13596 6237 6238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13595 7451 6238 6237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13594 7451 6238 6237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13593 6237 6238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13592 7451 7207 6239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13591 6302 6239 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13590 7451 6239 6302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13589 7451 6239 6302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13588 6302 6239 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13587 7451 7207 6171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13586 6172 6171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13585 7451 6171 6172 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13584 7451 6171 6172 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13583 6172 6171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13582 7451 7207 6244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13581 6243 6244 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13580 7451 6244 6243 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13579 7451 6244 6243 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13578 6243 6244 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13577 7451 7207 6245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13576 6528 6245 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13575 7451 6245 6528 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13574 7451 6245 6528 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13573 6528 6245 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13572 7451 7207 7134 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13571 7133 7134 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13570 7451 7134 7133 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13569 7451 7134 7133 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13568 7133 7134 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13567 7451 7207 7198 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13566 7197 7198 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13565 7451 7198 7197 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13564 7451 7198 7197 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13563 7197 7198 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13562 7451 7207 7200 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13561 7199 7200 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13560 7451 7200 7199 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13559 7451 7200 7199 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13558 7199 7200 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13557 4646 4979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13556 7451 6173 4645 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13555 7451 4912 4648 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13554 4647 4912 4646 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13553 4645 4648 4647 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13552 4644 4647 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13551 2453 3837 2410 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13550 2410 2454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13549 7451 4589 2453 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13548 2452 2453 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13547 4594 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13546 4594 4441 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13545 7451 4448 4594 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13544 7451 4446 4594 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13543 7221 7379 7220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13542 7220 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13541 7451 7489 7221 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13540 7219 7221 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13539 6638 6885 6580 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13538 6580 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13537 7451 7034 6580 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13536 6637 6638 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13535 6579 7032 6638 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13534 6580 7024 6579 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13533 6846 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13532 6846 4447 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13531 7451 4377 6846 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13530 7451 4376 6846 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13529 7451 7207 7140 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13528 7141 7140 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13527 7451 7140 7141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13526 7451 7140 7141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13525 7141 7140 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13524 7451 7207 7206 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13523 7205 7206 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13522 7451 7206 7205 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13521 7451 7206 7205 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13520 7205 7206 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13519 7451 7207 7209 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13518 7208 7209 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13517 7451 7209 7208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13516 7451 7209 7208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13515 7208 7209 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13514 7451 6739 4753 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13513 5280 4753 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13512 7451 4753 5280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13511 7451 4753 5280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13510 5280 4753 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13509 2157 2383 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13508 2157 2159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13507 7451 2514 2157 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13506 7451 2304 2157 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13505 7451 819 766 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13504 766 765 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13503 1022 1153 766 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13502 764 905 1022 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13501 766 1029 764 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13500 7451 6739 4767 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13499 5296 4767 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13498 7451 4767 5296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13497 7451 4767 5296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13496 5296 4767 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13495 7451 6739 6725 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13494 7194 6725 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13493 7451 6725 7194 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13492 7451 6725 7194 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13491 7194 6725 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13490 7451 6739 6740 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13489 7207 6740 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13488 7451 6740 7207 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13487 7451 6740 7207 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13486 7207 6740 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13485 5250 5718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13484 7451 6266 5250 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13483 5249 5250 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13482 6258 6259 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13481 7451 6473 6258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13480 6700 6258 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13479 5063 5066 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13478 5059 5067 5060 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13477 7451 6392 5059 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13476 5067 5068 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13475 7451 5594 5068 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13474 7451 5065 5066 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13473 5064 5067 5063 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13472 5062 5068 5064 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13471 7451 5061 5062 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13470 5061 5064 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13469 5060 5068 5061 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13468 7451 5060 6392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13467 6392 5060 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13466 6578 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13465 6631 7379 6578 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13464 7451 7454 6631 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13463 4478 4479 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13462 4472 4480 4474 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13461 7451 6025 4472 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13460 4480 4481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13459 7451 4638 4481 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13458 7451 4475 4479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13457 4477 4480 4478 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13456 4476 4481 4477 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13455 7451 4473 4476 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13454 4473 4477 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13453 4474 4481 4473 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13452 7451 4474 6025 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13451 6025 4474 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13450 7451 1051 1053 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13449 1053 1052 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13448 1053 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13447 7451 5173 1053 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13446 6332 1053 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13445 454 455 410 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13444 410 893 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13443 7451 641 454 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13442 554 454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13441 7451 6553 6552 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13440 6521 6628 6522 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13439 6522 6553 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13438 6522 6552 6521 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13437 7451 6551 6522 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13436 6551 6628 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13435 7451 3958 2564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13434 2565 3957 2932 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13433 2563 2587 2565 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13432 2564 6030 2563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13431 6641 7489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13430 6641 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13429 7451 6968 6641 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13428 7451 325 29 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13427 470 281 9 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13426 9 325 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13425 9 29 470 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13424 7451 27 9 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13423 27 281 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13422 6696 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13421 6696 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13420 7451 6968 6696 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13419 5236 5233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13418 7451 5234 5236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13417 5235 5236 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13416 2954 5690 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13415 2954 2174 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13414 7451 4158 2954 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13413 828 1342 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13412 828 514 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13411 7451 515 828 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13410 2614 2685 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13409 7451 2613 2614 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13408 2612 2614 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13407 3730 3729 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13406 7451 4732 3730 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13405 4264 3730 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13404 7451 7422 6684 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13403 6684 6683 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13402 7451 6882 6684 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13401 6682 6684 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13400 7451 7218 6563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13399 6563 6562 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13398 7451 6641 6563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13397 6598 6563 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13396 1342 1768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13395 7451 1435 1342 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13394 1826 2103 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13393 1826 2033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13392 7451 4081 1826 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13391 7451 7162 1826 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13390 1858 1257 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13389 7451 1258 1858 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13388 7451 899 145 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13387 461 900 116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13386 116 899 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13385 116 145 461 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13384 7451 146 116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13383 146 900 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13382 6259 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13381 6259 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13380 7451 5454 6259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13379 7451 6333 6259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13378 7451 793 531 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13377 721 531 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13376 7451 531 721 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13375 7451 531 721 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13374 721 531 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13373 7451 721 158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13372 4081 158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13371 7451 158 4081 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13370 7451 158 4081 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13369 4081 158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13368 7451 721 722 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13367 4600 722 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13366 7451 722 4600 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13365 7451 722 4600 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13364 4600 722 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13363 6673 6731 6675 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13362 6675 7034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13361 7451 7033 6675 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13360 6672 6673 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13359 6674 7032 6673 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13358 6675 6817 6674 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13357 3078 3077 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13356 7451 3483 3078 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13355 3137 3078 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13354 2812 2814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13353 7451 2811 2812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13352 3501 2812 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13351 7451 7387 7348 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13350 7348 7512 7356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13349 5859 6600 7033 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13348 5901 6047 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13347 7451 5901 5859 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13346 4496 4499 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13345 4492 4500 4493 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13344 7451 4782 4492 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13343 4500 4501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13342 7451 4561 4501 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13341 7451 4498 4499 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13340 4497 4500 4496 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13339 4495 4501 4497 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13338 7451 4494 4495 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13337 4494 4497 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13336 4493 4501 4494 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13335 7451 4493 4782 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13334 4782 4493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13333 151 470 117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13332 117 576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13331 7451 464 151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13330 126 151 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13329 7451 1572 1573 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13328 1573 2035 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13327 2958 7114 1573 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13326 1571 2174 2958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13325 1573 1837 1571 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13324 7451 2684 2331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13323 2331 2687 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13322 7451 4000 2331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13321 2328 2331 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13320 2928 5887 2927 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13319 3080 3226 2928 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13318 2928 3081 3080 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13317 2927 2926 2928 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13316 2927 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13315 7451 5274 2927 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13314 6443 7452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13313 7488 7489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13312 3992 4215 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13311 4067 4207 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13310 7463 7462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13309 1618 1976 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13308 7451 1049 1618 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13307 7451 2723 2100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13306 2100 2099 2101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13305 6271 6576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13304 7451 6652 6271 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13303 7451 6600 5824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13302 5827 6599 5826 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13301 5825 6406 5827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13300 5824 5832 5825 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13299 1112 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13298 7451 1908 1112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13297 1445 1112 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13296 7451 1111 1445 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13295 7451 5685 5383 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13294 5383 5467 5384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13293 5891 5384 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13292 4529 5216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13291 7451 6388 4530 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13290 7451 4912 4553 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13289 4552 4912 4529 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13288 4530 4553 4552 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13287 4635 4552 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13286 2988 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13285 7451 6333 2988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13284 4914 5055 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13283 7451 6392 4911 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13282 7451 4912 4915 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13281 4913 4912 4914 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13280 4911 4915 4913 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13279 5065 4913 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13278 2842 3484 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13277 7451 3483 2842 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13276 3912 4360 3914 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13275 3914 3913 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13274 7451 6326 3912 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13273 3911 3912 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13272 4370 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13271 4370 4603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13270 7451 4600 4370 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13269 7451 7114 4370 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13268 5363 5735 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13267 5708 5734 5363 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13266 7451 5876 5708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13265 5855 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13264 6384 6394 5855 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13263 7451 5882 6384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13262 796 1449 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13261 7451 4376 796 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13260 1384 796 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13259 7451 1034 705 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13258 3637 829 681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13257 681 1034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13256 681 705 3637 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13255 7451 703 681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13254 703 829 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13253 4507 4986 4508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13252 4508 6408 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13251 7451 6407 4508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13250 4998 4507 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13249 4506 4987 4507 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13248 4508 4984 4506 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13247 7451 4728 4731 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13246 4731 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13245 7451 7114 4731 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13244 6600 4731 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13243 6989 7387 6963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13242 6963 6990 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13241 7451 6992 6963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13240 7343 6989 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13239 6962 6991 6989 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13238 6963 7045 6962 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13237 7451 1304 812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13236 812 1906 872 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13235 1575 872 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13234 4785 5378 4815 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13233 4784 4783 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13232 7451 4784 4785 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13231 1978 2189 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13230 7451 2256 1978 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13229 2332 1978 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13228 4106 2602 2411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13227 2411 2457 4106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13226 7451 2456 2411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13225 604 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13224 7451 1908 604 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13223 728 604 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13222 7451 762 450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13221 1023 1068 409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13220 409 762 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13219 409 450 1023 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13218 7451 451 409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13217 451 1068 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13216 7451 1574 1439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13215 1439 1575 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13214 7451 2602 1439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13213 2040 1439 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13212 1622 1834 1592 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13211 1592 1620 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13210 7451 1619 1592 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13209 1974 1622 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13208 1591 5467 1622 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13207 1592 1618 1591 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13206 7451 2037 1836 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13205 1836 1835 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13204 1836 1896 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13203 7451 1899 1836 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13202 2333 1836 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13201 2671 2673 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13200 2665 2674 2668 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13199 7451 2664 2665 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13198 2674 2675 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13197 7451 2672 2675 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13196 7451 2669 2673 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13195 2670 2674 2671 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13194 2666 2675 2670 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13193 7451 2667 2666 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13192 2667 2670 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13191 2668 2675 2667 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13190 7451 2668 2664 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13189 2664 2668 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13188 302 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13187 319 372 302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13186 301 370 319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13185 7451 953 301 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13184 462 319 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13183 700 698 674 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13182 674 699 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13181 7451 1341 700 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13180 768 700 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13179 6547 6621 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13178 6541 6592 6616 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13177 7451 6617 6541 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13176 6592 6619 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13175 7451 6622 6619 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13174 7451 6620 6621 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13173 6590 6592 6547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13172 6548 6619 6590 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13171 7451 6589 6548 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13170 6589 6590 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13169 6616 6619 6589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13168 7451 6616 6617 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13167 6617 6616 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13166 5291 7511 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13165 5291 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13164 7451 5826 5291 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13163 3756 3771 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13162 3773 4697 3756 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13161 3755 4695 3773 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13160 7451 3770 3755 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13159 3769 3773 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13158 2560 6025 2559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13157 2583 3499 2560 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13156 2560 3135 2583 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13155 2559 2926 2560 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13154 2559 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13153 7451 5137 2559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13152 5676 5829 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13151 7451 5675 5676 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13150 1652 1203 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13149 7451 1569 1652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13148 7451 2082 2079 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13147 3159 2081 2083 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13146 2083 2082 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13145 2083 2079 3159 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13144 7451 2080 2083 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13143 2080 2081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13142 6240 6241 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13141 7451 6386 6240 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13140 6683 6240 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13139 3609 4838 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13138 3626 4413 3609 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13137 3608 4411 3626 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13136 7451 3978 3608 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13135 3625 3626 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13134 5374 5371 5375 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13133 5372 5818 5374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13132 5373 5819 5372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13131 7451 5815 5373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_13130 5679 5375 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13129 6248 6247 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13128 7451 6957 6248 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13127 6562 6248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13126 3704 4971 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13125 3703 4413 3704 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13124 3702 4411 3703 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13123 7451 3705 3702 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13122 3701 3703 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13121 1597 2602 1976 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13120 1661 2111 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13119 7451 1661 1597 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13118 7451 6266 4693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13117 4693 4828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13116 4732 7162 4693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13115 4692 4790 4732 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13114 4693 5016 4692 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13113 3166 4984 3123 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13112 3123 4987 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13111 7451 4986 3166 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13110 3326 3166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13109 6401 6399 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13108 7451 6531 6401 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13107 6400 6401 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13106 5684 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13105 5683 7383 5684 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13104 7451 7454 5683 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13103 3932 5134 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13102 3980 4413 3932 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13101 3931 4411 3980 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13100 7451 4112 3931 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13099 3979 3980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13098 6567 6568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13097 7451 6569 6567 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13096 6532 6567 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13095 6282 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13094 6328 7383 6282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13093 7451 6676 6328 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13092 5394 5470 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13091 5393 6058 5394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13090 7451 5693 5393 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13089 7451 6518 6374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13088 6372 6443 6373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13087 6373 6518 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13086 6373 6374 6372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13085 7451 6371 6373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13084 6371 6443 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13083 1039 2591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13082 7451 1577 1039 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13081 1355 1039 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13080 3990 4360 3940 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13079 3940 3992 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13078 7451 5307 3990 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13077 3989 3990 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_13076 934 1168 1385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13075 987 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13074 7451 987 934 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13073 3068 3066 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13072 7451 3067 3068 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13071 3074 3068 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13070 1058 1866 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13069 1079 1270 1058 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13068 1057 1341 1079 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13067 7451 1342 1057 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13066 1266 1079 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13065 2519 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13064 2520 2946 2519 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13063 7451 5137 2520 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13062 7451 1636 1635 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13061 1635 1633 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13060 7451 1634 1635 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13059 1598 1635 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13058 7451 1641 1640 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13057 1640 2008 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13056 7451 1855 1640 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13055 4987 1640 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13054 7451 5537 5538 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13053 5538 5751 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13052 7451 6955 5538 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13051 5539 5538 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13050 7217 7219 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13049 7218 7377 7217 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13048 7451 7420 7218 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13047 5916 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13046 7451 6061 5916 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_13045 7164 5916 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13044 6857 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13043 6885 7379 6857 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13042 7451 7481 6885 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13041 3429 3742 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13040 3733 3428 3429 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13039 7451 3427 3733 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13038 6285 6337 6339 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13037 6284 6338 6285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13036 7451 7334 6284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13035 4382 4407 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13034 4380 4409 4405 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13033 7451 4642 4380 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13032 4409 4408 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13031 7451 4488 4408 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_13030 7451 4765 4407 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13029 4395 4409 4382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13028 4381 4408 4395 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13027 7451 4394 4381 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13026 4394 4395 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13025 4405 4408 4394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13024 7451 4405 4642 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13023 4642 4405 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13022 3739 3993 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13021 3467 3466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13020 7451 3467 3468 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_13019 3465 3463 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13018 7451 3465 3449 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13017 3449 3468 3462 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13016 3462 3467 3448 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13015 3447 4148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13014 7451 3511 4148 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13013 4148 3511 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13012 3448 3460 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13011 3460 3462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13010 7451 7500 3460 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13009 3511 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_13008 3511 3468 3447 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13007 3460 3467 3511 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_13006 2872 3819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13005 5619 1304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13004 7287 6991 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13003 2544 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13002 2681 2541 2544 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13001 7451 2542 2681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_13000 41 162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12999 7451 3120 41 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12998 480 338 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12997 7451 2875 480 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12996 130 193 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12995 7451 2817 130 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12994 7451 6869 6818 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12993 6817 6965 6816 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12992 6816 6869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12991 6816 6818 6817 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12990 7451 6815 6816 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12989 6815 6965 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12988 6404 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12987 6570 6566 6404 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12986 7451 7453 6570 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12985 905 949 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12984 7451 951 905 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12983 5385 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12982 2541 1109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12981 7451 1111 2541 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12980 295 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12979 7451 3346 295 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12978 5729 6965 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12977 5729 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12976 7451 6968 5729 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12975 2472 2813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12974 7451 4934 2472 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12973 2688 2472 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12972 6890 7278 6860 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12971 6860 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12970 7451 7034 6860 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12969 6888 6890 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12968 6859 7032 6890 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12967 6860 7274 6859 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12966 463 464 414 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12965 414 512 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12964 7451 571 414 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12963 566 463 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12962 413 576 463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12961 414 470 413 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12960 949 1809 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12959 7451 1271 949 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12958 5858 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12957 5988 7383 5858 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12956 7451 7462 5988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12955 6253 7494 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12954 6253 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12953 7451 6980 6253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12952 1619 1501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12951 7451 1500 1619 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12950 5734 1489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12949 7451 1694 5734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12948 3389 3160 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12947 7451 3159 3389 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12946 169 4979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12945 7451 4934 168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12944 7451 6344 170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12943 188 6344 169 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12942 168 170 188 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12941 584 188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12940 677 4834 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12939 7451 4161 676 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12938 7451 6344 720 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12937 718 6344 677 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12936 676 720 718 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12935 785 718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12934 4238 6166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12933 4249 6165 4238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12932 7451 5069 4249 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12931 7451 1168 399 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12930 7451 1449 400 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12929 399 400 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12928 4518 4081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12927 7451 4437 4518 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12926 4819 5178 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12925 4819 4726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12924 7451 4724 4819 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12923 419 5274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12922 7451 1449 418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12921 7451 6344 474 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12920 473 6344 419 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12919 418 474 473 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12918 527 473 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12917 2001 5043 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12916 7451 2111 2000 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12915 7451 6344 2048 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12914 2047 6344 2001 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12913 2000 2048 2047 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12912 2118 2047 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12911 7251 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12910 7278 7379 7251 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12909 7451 7480 7278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12908 1356 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12907 1356 1041 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12906 7451 1040 1356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12905 7451 4589 1356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12904 1236 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12903 1236 2392 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12902 7451 1384 1236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12901 7451 2881 1236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12900 2978 4852 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12899 3002 4413 2978 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12898 2977 4411 3002 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12897 7451 3001 2977 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12896 3000 3002 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12895 2818 3348 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12894 7451 3343 2818 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12893 2817 2818 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12892 7451 6940 5802 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12891 5802 5801 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12890 7451 6158 5802 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12889 5952 5802 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12888 7451 7391 7115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12887 7115 7164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12886 7115 7113 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12885 7451 7114 7115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12884 7174 7115 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12883 2511 2926 2513 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12882 2513 3135 2512 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12881 2512 3500 2513 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12880 2511 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12879 7451 5055 2511 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12878 2513 6392 2511 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12877 2510 2512 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12876 7451 642 505 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12875 558 507 508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12874 508 642 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12873 508 505 558 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12872 7451 506 508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12871 506 507 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12870 1856 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12869 7451 1858 1856 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12868 1855 1856 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12867 1285 2095 1286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12866 1286 1287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12865 7451 1284 1285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12864 1489 1285 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12863 5398 5431 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12862 5396 5432 5425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12861 7451 5746 5396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12860 5432 5433 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12859 7451 5518 5433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12858 7451 5429 5431 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12857 5427 5432 5398 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12856 5397 5433 5427 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12855 7451 5426 5397 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12854 5426 5427 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12853 5425 5433 5426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12852 7451 5425 5746 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12851 5746 5425 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12850 3157 3722 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12849 7451 3321 3157 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12848 3156 3157 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12847 2535 2536 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12846 7451 2811 2535 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12845 3456 2535 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12844 3231 3989 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12843 7451 3502 3231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12842 3232 3231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12841 7451 4694 2014 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12840 2014 2524 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12839 7451 2228 2014 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12838 2139 2014 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12837 7451 2576 1863 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12836 1863 2416 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12835 7451 2220 1863 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12834 2647 1863 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12833 549 600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12832 547 599 593 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12831 7451 3820 547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12830 599 601 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12829 7451 598 601 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12828 7451 915 600 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12827 596 599 549 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12826 548 601 596 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12825 7451 595 548 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12824 595 596 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12823 593 601 595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12822 7451 593 3820 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12821 3820 593 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12820 7451 2733 2595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12819 2595 4367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12818 7451 4724 2595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12817 2592 2595 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12816 7451 2880 2393 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12815 2393 2392 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12814 2393 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12813 7451 2881 2393 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12812 2536 2393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12811 7451 1680 268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12810 1144 266 267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12809 267 1680 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12808 267 268 1144 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12807 7451 265 267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12806 265 266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12805 2996 4695 2976 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12804 2976 3481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12803 7451 3077 2996 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12802 3079 2996 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12801 7451 3814 1158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12800 1158 2174 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12799 1158 4158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12798 7451 5690 1158 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12797 1732 1158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12796 2324 2541 2272 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12795 2272 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12794 7451 2322 2324 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12793 3023 2324 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12792 7451 312 173 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12791 1465 1332 175 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12790 175 312 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12789 175 173 1465 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12788 7451 174 175 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12787 174 1332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12786 3252 3655 3251 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12785 3251 4569 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12784 7451 3659 3252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12783 3348 3252 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12782 4636 4637 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12781 4631 4639 4630 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12780 7451 6388 4631 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12779 4639 4640 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12778 7451 4638 4640 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12777 7451 4635 4637 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12776 4633 4639 4636 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12775 4634 4640 4633 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12774 7451 4632 4634 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12773 4632 4633 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12772 4630 4640 4632 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12771 7451 4630 6388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12770 6388 4630 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12769 4924 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12768 4923 5273 4924 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12767 7451 6173 4923 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12766 6103 6169 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12765 6761 6168 6103 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12764 7451 6125 6761 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12763 5379 5377 5381 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12762 5380 6910 5379 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12761 7451 5378 5380 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12760 6863 6991 6915 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12759 6864 7512 6863 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12758 7451 7387 6864 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12757 6914 6915 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12756 3110 3109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12755 7451 4852 3112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12754 7451 3667 3113 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12753 3111 3667 3110 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12752 3112 3113 3111 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12751 3108 3111 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12750 2258 5467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12749 2457 2256 2258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12748 7451 2257 2457 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12747 7451 7471 7472 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12746 7470 7473 7446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12745 7446 7471 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12744 7446 7472 7470 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12743 7451 7467 7446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12742 7467 7473 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12741 5897 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12740 5897 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12739 7451 6980 5897 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12738 5315 5840 5263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12737 5263 7108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12736 7451 5842 5263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12735 5876 5315 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12734 5262 5841 5315 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12733 5263 6133 5262 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12732 7102 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12731 7101 7428 7102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12730 7451 7493 7101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12729 75 2134 181 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12728 76 3546 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12727 7451 76 75 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12726 1893 2813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12725 7451 2536 1893 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12724 6194 7114 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12723 6194 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12722 7451 6266 6194 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12721 4853 5369 4797 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12720 4797 4852 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12719 7451 5226 4853 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12718 5967 4853 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12717 4675 4673 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12716 7451 4674 4675 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12715 6405 4675 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12714 4564 4986 4535 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12713 4535 4566 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12712 7451 5085 4535 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12711 4809 4564 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12710 4534 4987 4564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12709 4535 4984 4534 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12708 3440 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12707 3502 4669 3440 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12706 7451 3500 3502 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12705 3279 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12704 3322 4669 3279 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12703 7451 3645 3322 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12702 5694 6773 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12701 7451 6056 5694 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12700 5693 5694 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12699 7451 1700 1590 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12698 1590 1968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12697 1750 1967 1590 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12696 1589 5735 1750 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12695 1590 5734 1589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12694 2826 3214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12693 2841 3212 2826 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12692 7451 6617 2841 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12691 7451 3352 3115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12690 3115 4158 3114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12689 3428 3114 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12688 2257 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12687 2257 2591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12686 7451 2880 2257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12685 7451 2881 2257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12684 1734 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12683 7451 1732 1734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12682 1733 1734 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12681 3039 3119 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12680 7451 3266 3039 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12679 3037 3039 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12678 2506 2502 2503 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12677 3407 2504 2506 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12676 2506 2505 3407 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12675 2503 3138 2506 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12674 2503 2789 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12673 7451 2794 2503 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12672 2380 2986 2507 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12671 2379 2520 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12670 7451 2379 2380 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12669 6571 6572 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12668 7451 6570 6571 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12667 6644 6571 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12666 4668 5093 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12665 7451 4732 4668 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12664 4667 4668 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12663 7451 6979 6978 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12662 6978 6980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12661 7451 7475 6978 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12660 6954 6978 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12659 7451 7234 6709 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12658 6709 6707 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12657 7451 6708 6709 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12656 6902 6709 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12655 7451 7283 7284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12654 7427 7284 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12653 7451 7284 7427 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12652 7451 7284 7427 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12651 7427 7284 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12650 7451 7427 7429 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12649 7428 7429 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12648 7451 7429 7428 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12647 7451 7429 7428 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12646 7428 7429 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12645 7451 7427 7380 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12644 7379 7380 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12643 7451 7380 7379 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12642 7451 7380 7379 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12641 7379 7380 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12640 7451 1764 1722 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12639 1722 1765 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12638 3178 7114 1722 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12637 1721 2174 3178 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12636 1722 1837 1721 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12635 772 1187 773 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12634 773 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12633 7451 771 772 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12632 824 772 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12631 1208 1501 1176 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12630 1176 1365 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12629 7451 1500 1208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12628 2179 1208 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12627 7451 1954 1955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12626 6166 1952 1953 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12625 1953 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12624 1953 1955 6166 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12623 7451 1951 1953 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12622 1951 1952 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12621 4061 4062 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12620 4055 4063 4057 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12619 7451 4069 4055 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12618 4063 4064 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12617 7451 4561 4064 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12616 7451 4059 4062 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12615 4060 4063 4061 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12614 4056 4064 4060 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12613 7451 4058 4056 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12612 4058 4060 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12611 4057 4064 4058 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12610 7451 4057 4069 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12609 4069 4057 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12608 6105 6393 6967 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12607 6104 6315 6105 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12606 7451 6394 6104 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12605 4988 4986 4947 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12604 4947 4985 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12603 7451 5085 4947 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12602 5879 4988 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12601 4946 4987 4988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12600 4947 4984 4946 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12599 3443 3506 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12598 3441 3507 3504 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12597 7451 3727 3441 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12596 3507 3508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12595 7451 3581 3508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12594 7451 3648 3506 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12593 3455 3507 3443 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12592 3442 3508 3455 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12591 7451 3453 3442 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12590 3453 3455 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12589 3504 3508 3453 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12588 7451 3504 3727 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12587 3727 3504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12586 7097 7144 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12585 7098 7372 7097 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12584 7451 7420 7098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12583 2881 2111 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12582 4000 2686 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12581 3742 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12580 1271 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12579 7451 3814 1271 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12578 5917 6061 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12577 5467 7162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12576 6017 7335 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12575 6017 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12574 7451 6968 6017 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12573 2743 4934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12572 2743 5994 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12571 7451 6133 2743 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12570 6122 6380 6098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12569 6098 7034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12568 7451 7033 6098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12567 6096 6122 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12566 6097 7032 6122 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12565 6098 6521 6097 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12564 6431 6474 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12563 6476 6894 6431 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12562 7451 6901 6476 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12561 4509 4726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12560 7451 4724 4509 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12559 4582 4509 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12558 471 1085 417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12557 417 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12556 7451 831 471 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12555 654 471 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12554 7451 4158 1327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12553 1327 3427 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12552 1373 1371 1327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12551 1326 5467 1373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12550 1327 1372 1326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12549 1040 963 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12548 1040 1292 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12547 7451 4081 1040 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12546 7451 5841 1040 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12545 1584 3135 1642 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12544 1583 1959 1584 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12543 7451 1736 1583 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12542 1684 1642 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12541 7451 2932 2933 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12540 2933 3636 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12539 7451 3637 2933 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12538 2999 2933 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12537 380 1085 381 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12536 381 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12535 7451 775 380 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12534 469 380 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12533 7312 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12532 7311 7379 7312 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12531 7451 7475 7311 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12530 2084 2140 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12529 7451 2085 2084 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12528 2217 2084 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12527 2742 2739 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12526 7451 2738 2742 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12525 2741 2742 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12524 7451 2602 2338 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12523 7451 4161 2194 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12522 2338 2194 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12521 5470 7388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12520 3500 4861 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12519 3644 4716 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12518 7451 1029 694 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12517 694 1145 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12516 7451 829 694 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12515 691 694 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12514 6702 6841 6703 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12513 6701 6700 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12512 7451 6701 6702 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12511 7451 6980 2107 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12510 2107 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12509 2319 2322 2107 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12508 2106 2543 2319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12507 2107 2541 2106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12506 3499 4502 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12505 2949 4504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12504 6809 6812 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12503 6805 6813 6806 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12502 7451 6804 6805 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12501 6813 6814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12500 7451 7189 6814 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12499 7451 6811 6812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12498 6810 6813 6809 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12497 6808 6814 6810 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12496 7451 6807 6808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12495 6807 6810 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12494 6806 6814 6807 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12493 7451 6806 6804 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12492 6804 6806 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12491 6123 6124 6101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12490 6101 7034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12489 7451 7033 6101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12488 6099 6123 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12487 6100 7032 6123 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12486 6101 6678 6100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12485 284 653 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12484 283 654 284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12483 7451 777 283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12482 7451 5691 5692 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12481 5692 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12480 7451 5690 5692 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12479 6337 5692 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12478 2924 6388 2923 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12477 2922 3644 2924 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12476 2924 3135 2922 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12475 2923 2926 2924 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12474 2923 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12473 7451 5216 2923 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12472 2885 2951 2835 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12471 2835 6342 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12470 7451 2884 2885 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12469 2887 2885 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12468 4755 4959 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12467 4755 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12466 7451 5826 4755 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12465 5895 6107 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12464 7451 6180 5895 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12463 5400 5435 5436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12462 5401 5818 5400 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12461 5399 5819 5401 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12460 7451 5815 5399 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_12459 5434 5436 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12458 1727 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12457 7451 3646 1727 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12456 4843 5369 4796 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12455 4796 4841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12454 7451 5226 4843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12453 5413 4843 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12452 5077 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12451 5234 5273 5077 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12450 7451 5882 5234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12449 1474 1550 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12448 1474 1473 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12447 7451 1686 1474 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12446 3347 5225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12445 3347 3917 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12444 7451 3170 3347 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12443 519 654 520 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12442 520 653 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12441 7451 833 519 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12440 706 519 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12439 7451 4368 4357 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12438 4357 5085 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12437 4357 4367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12436 7451 4985 4357 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12435 4401 4357 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12434 1447 1445 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12433 1448 2179 1447 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12432 1446 2541 1448 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12431 7451 2543 1446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12430 1444 1448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12429 204 237 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12428 202 236 230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12427 7451 1304 202 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12426 236 238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12425 7451 669 238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12424 7451 233 237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12423 235 236 204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12422 203 238 235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12421 7451 231 203 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12420 231 235 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12419 230 238 231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12418 7451 230 1304 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12417 1304 230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12416 2278 2661 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12415 2429 2658 2278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12414 7451 2502 2429 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12413 7451 3769 2422 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12412 2422 2507 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12411 7451 2508 2422 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12410 3549 2422 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12409 2869 2813 2815 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12408 2815 2814 2869 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12407 7451 2872 2815 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12406 5983 5984 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12405 7451 6253 5983 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12404 5982 5983 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12403 5390 6845 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12402 5389 5387 5390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12401 5388 6846 5389 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12400 7451 5385 5388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12399 5386 5389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12398 7451 5681 5682 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12397 5682 5683 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12396 7451 6185 5682 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12395 5810 5682 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12394 5614 5616 5570 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12393 5570 5617 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12392 7451 5889 5614 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12391 6893 5614 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12390 2930 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12389 3483 2929 2930 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12388 7451 5887 3483 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12387 6000 6014 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12386 6015 6375 6000 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12385 7451 7420 6015 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12384 7451 1574 1576 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12383 1576 1575 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12382 7451 2255 1576 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12381 2042 1576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12380 3597 3734 3599 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12379 3599 3733 3598 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12378 3598 3732 3599 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12377 3597 3920 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12376 7451 4077 3597 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12375 3599 3967 3597 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12374 6980 3598 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12373 7451 1736 176 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12372 1332 1413 178 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12371 178 1736 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12370 178 176 1332 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12369 7451 177 178 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12368 177 1413 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12367 4800 4858 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12366 4798 4859 4855 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12365 7451 5160 4798 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12364 4859 4860 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12363 7451 5531 4860 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12362 7451 4857 4858 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12361 4813 4859 4800 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12360 4799 4860 4813 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12359 7451 4812 4799 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12358 4812 4813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12357 4855 4860 4812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12356 7451 4855 5160 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12355 5160 4855 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12354 5189 5554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12353 7451 5189 5188 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12352 5187 5331 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12351 7451 5187 5115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12350 5115 5188 5185 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12349 5185 5189 5114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12348 5113 7390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12347 7451 5181 7390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12346 7390 5181 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12345 5114 5182 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12344 5182 5185 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12343 7451 7500 5182 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12342 5181 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12341 5181 5188 5113 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12340 5182 5189 5181 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12339 5701 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12338 5751 7383 5701 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12337 7451 6628 5751 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12336 6113 6538 6114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12335 6134 6533 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12334 7451 6134 6113 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12333 2284 2602 2813 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12332 2340 4161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12331 7451 2340 2284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12330 2009 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12329 7451 1858 2009 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12328 2094 2093 4986 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12327 2092 2090 2094 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12326 7451 2091 2092 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12325 7451 181 22 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12324 900 272 7 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12323 7 181 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12322 7 22 900 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12321 7451 19 7 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12320 19 272 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12319 6533 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12318 7451 7384 6533 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12317 2834 2953 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12316 2866 2865 2834 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12315 7451 3108 2866 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12314 1749 3159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12313 1749 3160 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12312 7451 1567 1749 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12311 7451 3179 2955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12310 2955 2954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12309 7451 2995 2955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12308 2953 2955 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12307 6907 5718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12306 7451 6133 6907 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12305 4367 7108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12304 4367 4603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12303 7451 4600 4367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12302 5256 5834 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12301 7451 4998 5256 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12300 5807 6628 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12299 5807 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12298 7451 6968 5807 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12297 7451 7212 6313 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12296 6313 6310 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12295 7451 6831 6313 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12294 6309 6313 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12293 7451 6948 6636 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12292 6636 6633 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12291 7451 6741 6636 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12290 6632 6636 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12289 4772 4771 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12288 7451 4923 4772 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12287 5079 4772 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12286 1235 1236 1177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12285 7451 1440 1177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12284 1177 1441 1235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12283 6407 1235 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12282 7229 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12281 7430 7228 7229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12280 7451 7489 7430 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12279 6196 6195 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12278 7451 6194 6196 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12277 6193 6196 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12276 7451 6322 5980 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12275 5980 6037 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12274 7451 6391 5980 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12273 6032 5980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12272 7451 5757 5253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12271 5253 5252 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12270 7451 5386 5253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12269 5251 5253 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12268 1851 1435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12267 1851 1968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12266 7451 1700 1851 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12265 7451 1688 1851 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12264 1701 4726 1702 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12263 1702 2103 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12262 7451 4773 1701 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12261 1700 1701 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12260 4597 1915 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12259 4597 1775 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12258 7451 4446 4597 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12257 7451 3742 4597 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12256 7451 571 308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12255 308 512 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12254 823 464 308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12253 307 576 823 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12252 308 470 307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12251 542 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12250 568 1187 542 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12249 7451 771 568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12248 5608 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12247 5608 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12246 7451 5160 5608 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12245 7451 6333 5608 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12244 6913 6912 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12243 7451 7168 6913 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12242 6910 6913 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12241 6411 6652 6990 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12240 6412 6410 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12239 7451 6412 6411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12238 3489 3562 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12237 7451 3563 3489 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12236 3487 3489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12235 2950 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12234 3238 4669 2950 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12233 7451 3646 3238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12232 1960 2424 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12231 7451 2133 1960 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12230 1959 1960 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12229 5975 5977 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12228 5970 5979 5971 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12227 7451 5969 5970 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12226 5979 5978 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12225 7451 6693 5978 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12224 7451 5974 5977 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12223 5976 5979 5975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12222 5973 5978 5976 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12221 7451 5972 5973 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12220 5972 5976 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12219 5971 5978 5972 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12218 7451 5971 5969 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12217 5969 5971 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12216 2864 3233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12215 7451 2861 2864 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12214 2862 2864 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12213 916 1976 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12212 7451 1049 916 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12211 1628 916 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12210 7451 558 559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12209 3632 554 541 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12208 541 558 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12207 541 559 3632 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12206 7451 556 541 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12205 556 554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12204 636 1728 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12203 1634 937 636 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12202 7451 1681 1634 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12201 1220 1257 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12200 7451 1258 1220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12199 1952 1220 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12198 7246 7261 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12197 7263 7411 7246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12196 7451 7420 7263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12195 6858 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12194 6886 7428 6858 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12193 7451 7466 6886 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12192 4144 4360 4097 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12191 4097 4143 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12190 7451 6646 4144 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12189 4142 4144 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12188 7451 5718 4229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12187 4229 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12186 7451 4934 4229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12185 4228 4229 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12184 1776 1775 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12183 7451 4446 1776 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12182 1911 1776 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12181 89 90 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12180 85 91 84 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12179 7451 286 85 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12178 91 92 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12177 7451 598 92 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12176 7451 656 90 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12175 87 91 89 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12174 88 92 87 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12173 7451 86 88 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12172 86 87 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12171 84 92 86 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12170 7451 84 286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12169 286 84 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12168 7451 5172 4867 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12167 4867 5171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12166 7451 5173 4867 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12165 5840 4867 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12164 4871 5695 4808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12163 4808 5470 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12162 7451 6344 4871 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12161 4869 4871 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12160 2391 2537 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12159 2956 2390 2391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12158 7451 7162 2956 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12157 7451 1852 65 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12156 1681 262 64 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12155 64 1852 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12154 64 65 1681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12153 7451 63 64 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12152 63 262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12151 3354 4673 3283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12150 3283 3352 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12149 7451 4148 3354 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12148 3351 3354 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12147 1305 1765 1306 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12146 1306 1579 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12145 7451 1304 1305 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12144 1508 1305 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12143 4363 4360 4362 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12142 4362 4361 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12141 7451 6469 4363 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12140 4359 4363 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12139 4589 6979 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12138 7451 6980 4589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12137 5617 5457 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12136 7451 6333 5617 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12135 680 696 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12134 1029 767 680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12133 7451 695 1029 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12132 3563 3142 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12131 7451 3143 3563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12130 909 776 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12129 909 777 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12128 7451 778 909 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12127 3870 3633 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12126 7451 3632 3870 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12125 6112 7114 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12124 6112 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12123 7451 6133 6112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12122 6147 6342 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12121 6988 6340 6147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12120 7451 6713 6988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12119 5286 7495 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12118 5286 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12117 7451 5826 5286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12116 7451 5235 5152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12115 5152 6451 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12114 7451 5434 5152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12113 5230 5152 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12112 2502 1826 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12111 2502 1825 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12110 7451 2315 2502 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12109 7451 1684 1685 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12108 1685 1813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12107 1682 1679 1685 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12106 1683 1680 1682 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12105 1685 1681 1683 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12104 6406 6768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12103 6406 6405 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12102 7451 6843 6406 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12101 7451 6907 6406 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12100 1956 2926 1958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12099 1958 3135 1957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12098 1957 3646 1958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12097 1956 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12096 7451 4834 1956 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12095 1958 6175 1956 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12094 2222 1957 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12093 7451 5837 5838 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12092 5838 6407 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12091 7451 6408 5838 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12090 6048 5838 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12089 1086 2853 1059 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12088 1059 2435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12087 7451 2133 1086 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12086 1085 1086 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12085 7451 3625 800 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12084 800 2290 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12083 1334 3546 800 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12082 799 3549 1334 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12081 800 1866 799 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12080 2682 2681 2683 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12079 2683 5467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12078 7451 2743 2682 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12077 3029 2682 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12076 3909 4277 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12075 7451 3909 3910 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12074 3908 3905 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12073 7451 3908 3906 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12072 3906 3910 3907 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12071 3907 3909 3904 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12070 3901 4718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12069 7451 3902 4718 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12068 4718 3902 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12067 3904 3903 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12066 3903 3907 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12065 7451 5100 3903 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12064 3902 5100 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12063 3902 3910 3901 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12062 3903 3909 3902 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_12061 3745 3744 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12060 3743 5000 3745 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12059 7451 4378 3743 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12058 7145 7428 7119 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12057 7119 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12056 7451 7480 7145 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12055 7144 7145 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12054 2376 2926 2378 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12053 2378 3135 2377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12052 2377 3645 2378 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12051 2376 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12050 7451 5043 2376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12049 2378 6035 2376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12048 2433 2377 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12047 2110 2813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12046 7451 2536 2110 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12045 2109 2110 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12044 611 4728 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12043 7451 5001 611 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12042 609 611 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12041 4676 5385 4677 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12040 4677 5619 4676 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12039 7451 6846 4677 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12038 7451 2241 1824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12037 1824 2101 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12036 7451 2165 1824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_12035 1823 1824 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12034 7451 7413 7409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12033 7411 7463 7412 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12032 7412 7413 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12031 7412 7409 7411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12030 7451 7410 7412 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12029 7410 7463 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_12028 4093 4130 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12027 4091 4132 4124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12026 7451 4207 4091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12025 4132 4131 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12024 7451 4561 4131 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_12023 7451 4206 4130 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12022 4128 4132 4093 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12021 4092 4131 4128 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12020 7451 4126 4092 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12019 4126 4128 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12018 4124 4131 4126 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_12017 7451 4124 4207 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12016 4207 4124 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12015 7451 3004 1715 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12014 1715 1740 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12013 1741 3546 1715 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12012 1714 1823 1741 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12011 1715 1866 1714 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12010 1432 1823 1433 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12009 1433 2023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12008 7451 1431 1432 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12007 1747 1432 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12006 4065 4360 4068 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12005 4068 4067 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12004 7451 5982 4065 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12003 4066 4065 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_12002 5854 6030 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12001 5877 6029 5854 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_12000 7451 5876 5877 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11999 2972 2686 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11998 2972 2688 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11997 7451 2687 2972 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11996 5501 5500 5502 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11995 5499 5498 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11994 7451 5499 5501 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11993 7451 7474 7272 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11992 7270 7424 7249 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11991 7249 7474 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11990 7249 7272 7270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11989 7451 7268 7249 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11988 7268 7424 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11987 7451 4679 4523 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11986 4525 4676 4524 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11985 4522 4604 4525 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11984 4523 4790 4522 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11983 4918 5369 4917 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11982 4917 4916 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11981 7451 5226 4918 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11980 5662 4918 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11979 7342 7508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11978 7451 7342 7341 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11977 7340 7343 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11976 7451 7340 7322 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11975 7322 7341 7339 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11974 7339 7342 7323 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11973 7321 7387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11972 7451 7337 7387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11971 7387 7337 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11970 7323 7338 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11969 7338 7339 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11968 7451 7500 7338 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11967 7337 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11966 7337 7341 7321 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11965 7338 7342 7337 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11964 281 2016 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11963 7451 3546 281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11962 6145 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11961 6181 6566 6145 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11960 7451 7462 6181 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11959 2707 2795 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11958 2707 2708 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11957 7451 2705 2707 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11956 6102 6676 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11955 6102 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11954 7451 6968 6102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11953 642 951 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11952 642 1029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11951 7451 1732 642 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11950 682 731 730 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11949 683 728 682 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11948 7451 729 683 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11947 790 730 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11946 7451 942 679 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11945 679 939 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11944 1680 685 679 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11943 678 1021 1680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11942 679 1022 678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11941 5083 5043 4930 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11940 4930 5832 5083 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11939 7451 4929 4930 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11938 7451 4600 4152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11937 4152 4603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11936 4152 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11935 7451 7114 4152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11934 5832 4152 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11933 155 654 118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11932 118 653 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11931 7451 777 155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11930 468 155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11929 7451 1565 1566 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11928 1566 1883 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11927 7451 1699 1566 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11926 1695 1566 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11925 7451 7460 7132 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11924 7129 7454 7116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11923 7116 7460 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11922 7116 7132 7129 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11921 7451 7128 7116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11920 7128 7454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11919 5018 5691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11918 7451 5841 5018 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11917 5016 5018 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11916 2326 2454 2273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11915 2273 5467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11914 7451 2325 2326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11913 2730 2326 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11912 1697 2164 1698 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11911 1698 1823 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11910 7451 2023 1698 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11909 1694 1697 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11908 1696 1695 1697 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11907 1698 1819 1696 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11906 114 142 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11905 112 124 141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11904 7451 3868 112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11903 124 125 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11902 7451 368 125 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11901 7451 3876 142 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11900 121 124 114 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11899 113 125 121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11898 7451 120 113 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11897 120 121 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11896 141 125 120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11895 7451 141 3868 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11894 3868 141 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11893 2945 2676 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11892 7451 2956 2945 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11891 6119 5659 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11890 7451 5655 6119 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11889 4579 4726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11888 7451 4724 4579 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11887 3615 3649 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11886 7451 3727 3614 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11885 7451 4577 3652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11884 3650 4577 3615 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11883 3614 3652 3650 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11882 3648 3650 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11881 4336 5127 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11880 7451 4782 4335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11879 7451 4577 4337 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11878 4356 4577 4336 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11877 4335 4337 4356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11876 4498 4356 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11875 3759 3804 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11874 7451 4069 3760 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11873 7451 4577 3805 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11872 3803 4577 3759 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11871 3760 3805 3803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11870 4059 3803 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11869 3967 4079 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11868 7451 3966 3967 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11867 4516 5385 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11866 5377 4594 4516 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11865 4515 4593 5377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11864 7451 6846 4515 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11863 5870 5805 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11862 7451 5708 5870 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11861 4209 4211 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11860 7451 4207 4208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11859 7451 4577 4212 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11858 4210 4577 4209 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11857 4208 4212 4210 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11856 4206 4210 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11855 3837 4934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11854 7451 4158 3837 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11853 4685 4698 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11852 4699 4697 4685 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11851 4684 4695 4699 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11850 7451 4696 4684 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11849 4694 4699 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11848 2568 3389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11847 7451 2596 2567 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11846 7451 5128 2601 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11845 2600 5128 2568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11844 2567 2601 2600 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11843 2597 2600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11842 3239 4070 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11841 7451 3238 3239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11840 6576 7162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11839 6576 7164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11838 7451 7391 6576 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11837 7112 7113 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11836 7505 7163 7112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11835 7451 7111 7505 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11834 7019 7311 6997 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11833 6997 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11832 7451 7034 6997 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11831 7018 7019 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11830 6996 7032 7019 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11829 6997 7366 6996 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11828 481 4376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11827 481 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11826 7451 3352 481 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11825 460 511 412 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11824 412 462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11823 7451 1032 412 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11822 695 460 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11821 411 1466 460 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11820 412 461 411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11819 5387 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11818 5387 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11817 7451 4447 5387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11816 7451 4934 5387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11815 1024 1021 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11814 1025 1022 1024 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11813 7451 1023 1025 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11812 3956 4488 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11811 7451 3956 3955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11810 3954 3953 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11809 7451 3954 3935 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11808 3935 3955 3951 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11807 3951 3956 3934 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11806 3933 4431 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11805 7451 3982 4431 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11804 4431 3982 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11803 3934 3949 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11802 3949 3951 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11801 7451 7500 3949 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11800 3982 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11799 3982 3955 3933 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11798 3949 3956 3982 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11797 5856 5884 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11796 6464 5885 5856 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11795 7451 6315 6464 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11794 7451 4934 4079 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11793 7451 4158 4080 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11792 4079 4080 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11791 1359 1577 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11790 7451 5000 1359 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11789 2789 1359 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11788 98 99 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11787 94 100 93 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11786 7451 190 94 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11785 100 101 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11784 7451 669 101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11783 7451 130 99 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11782 96 100 98 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11781 97 101 96 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11780 7451 95 97 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11779 95 96 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11778 93 101 95 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11777 7451 93 190 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11776 190 93 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11775 3010 3720 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11774 7451 3009 3010 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11773 3077 3010 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11772 1434 1568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11771 7451 1569 1434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11770 3212 1434 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11769 1545 3546 1546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11768 1546 1727 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11767 7451 3979 1546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11766 1543 1545 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11765 1544 2139 1545 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11764 1546 1866 1544 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11763 5609 5608 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11762 7451 6042 5609 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11761 6039 5609 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11760 4948 4991 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11759 5153 5381 4948 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11758 7451 6957 5153 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11757 3341 3466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11756 7451 3341 3342 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11755 3340 3338 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11754 7451 3340 3275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11753 3275 3342 3337 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11752 3337 3341 3274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11751 3273 4156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11750 7451 3334 4156 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11749 4156 3334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11748 3274 3335 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11747 3335 3337 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11746 7451 5100 3335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11745 3334 5100 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11744 3334 3342 3273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11743 3335 3341 3334 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11742 6949 6969 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11741 6948 7092 6949 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11740 7451 7420 6948 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11739 7451 1341 911 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11738 911 910 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11737 7451 909 911 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11736 3958 911 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11735 7159 7353 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11734 7451 7384 7159 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11733 7228 7159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11732 3117 3655 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11731 3463 3116 3117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11730 7451 3183 3463 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11729 4927 4834 4691 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11728 4691 5832 4927 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11727 7451 4722 4691 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11726 2231 2658 2230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11725 2230 2661 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11724 7451 2510 2231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11723 2229 2231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11722 1503 2541 1454 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11721 1454 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11720 7451 1628 1503 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11719 2174 1503 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11718 7451 3997 3944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11717 3944 4228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11716 5537 4156 3944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11715 3943 4149 5537 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11714 3944 5909 3943 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11713 7451 2880 2459 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11712 2459 2591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11711 2459 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11710 7451 2881 2459 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11709 2814 2459 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11708 1705 2541 1704 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11707 1704 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11706 7451 2035 1705 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11705 1880 1705 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11704 7451 7486 7487 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11703 7484 7489 7447 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11702 7447 7486 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11701 7447 7487 7484 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11700 7451 7482 7447 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11699 7482 7489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11698 2164 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11697 7451 2392 2164 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11696 7319 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11695 7320 7383 7319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11694 7451 7335 7320 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11693 1337 1422 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11692 7451 1474 1337 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11691 2558 2647 3411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11690 2557 2648 2558 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11689 7451 2655 2557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11688 6379 6625 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11687 6378 6942 6379 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11686 7451 7420 6378 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11685 3835 4305 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11684 7451 3835 3834 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11683 3833 3830 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11682 7451 3833 3754 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11681 3754 3834 3831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11680 3831 3835 3753 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11679 3752 3993 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11678 7451 3827 3993 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11677 3993 3827 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11676 3753 3828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11675 3828 3831 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11674 7451 7500 3828 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11673 3827 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11672 3827 3834 3752 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11671 3828 3835 3827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11670 6612 6611 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11669 7451 6612 6610 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11668 6609 6608 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11667 7451 6609 6574 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11666 6574 6610 6606 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11665 6606 6612 6573 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11664 6586 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11663 7451 6651 6652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11662 6652 6651 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11661 6573 6603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11660 6603 6606 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11659 7451 7500 6603 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11658 6651 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11657 6651 6610 6586 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11656 6603 6612 6651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11655 3184 3179 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11654 3184 3181 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11653 7451 3178 3184 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11652 6002 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11651 6241 6394 6002 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11650 7451 6025 6241 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11649 847 875 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11648 847 1632 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11647 7451 1114 847 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11646 893 829 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11645 893 1029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11644 7451 1145 893 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11643 1425 1682 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11642 1426 1479 1425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11641 7451 1556 1426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11640 2397 2398 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11639 2465 2813 2397 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11638 7451 2536 2465 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11637 5700 6600 5745 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11636 5699 6599 5700 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11635 5698 6406 5699 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11634 7451 5832 5698 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11633 5818 5745 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11632 3179 7114 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11631 3179 2816 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11630 7451 3023 3179 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11629 7451 7164 5120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11628 5120 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11627 5418 5138 5120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11626 5119 5275 5418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11625 5120 5273 5119 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11624 2171 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11623 2171 1970 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11622 7451 2033 2171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11621 7451 6333 2171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11620 6125 6407 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11619 7451 6408 6125 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11618 6707 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11617 6707 5718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11616 7451 4782 6707 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11615 7451 4934 6707 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11614 5991 6704 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11613 7451 6027 5991 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11612 4778 6894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11611 4779 4777 4778 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11610 7451 5242 4779 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11609 2562 6392 2561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11608 2708 3500 2562 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11607 2562 3135 2708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11606 2561 2926 2562 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11605 2561 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11604 7451 5055 2561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11603 7349 7390 7391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11602 7389 7388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11601 7451 7389 7349 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11600 1917 1915 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11599 7451 3742 1917 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11598 1914 1917 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11597 7451 894 891 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11596 6316 893 895 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11595 895 894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11594 895 891 6316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11593 7451 892 895 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11592 892 893 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11591 7426 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11590 7451 7494 7426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11589 7486 7426 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11588 7451 7164 6564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11587 6564 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11586 7451 7113 6564 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11585 6529 6564 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11584 5123 7388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11583 5178 7390 5123 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11582 7451 7384 5178 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11581 4828 4789 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11580 4828 5387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11579 7451 5620 4828 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11578 2500 4695 2501 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11577 2501 3129 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11576 7451 2841 2500 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11575 2785 2500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11574 7051 7236 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11573 7451 7287 7051 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11572 7049 7051 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11571 2104 2602 2105 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11570 2105 2536 2104 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11569 7451 2103 2105 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11568 2105 2814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11567 2370 2418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11566 7451 2504 2370 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11565 3071 2370 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11564 5530 5529 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11563 5525 5532 5524 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11562 7451 5523 5525 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11561 5532 5533 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11560 7451 5531 5533 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11559 7451 5676 5529 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11558 5528 5532 5530 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11557 5527 5533 5528 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11556 7451 5526 5527 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11555 5526 5528 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11554 5524 5533 5526 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11553 7451 5524 5523 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11552 5523 5524 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11551 6766 7109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11550 7451 7108 6766 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11549 7227 6766 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11548 5358 5360 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11547 5354 5361 5355 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11546 7451 7495 5354 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11545 5361 5362 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11544 7451 5594 5362 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11543 7451 5423 5360 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11542 5359 5361 5358 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11541 5357 5362 5359 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11540 7451 5356 5357 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11539 5356 5359 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11538 5355 5362 5356 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11537 7451 5355 7495 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11536 7495 5355 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11535 5623 6344 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11534 7111 1115 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11533 822 902 803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11532 803 1768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11531 7451 1435 803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11530 819 822 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11529 802 899 822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11528 803 900 802 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11527 6403 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11526 6402 6566 6403 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11525 7451 6628 6402 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11524 664 668 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11523 661 667 662 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11522 7451 1168 661 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11521 667 670 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11520 7451 669 670 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11519 7451 841 668 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11518 665 667 664 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11517 666 670 665 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11516 7451 663 666 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11515 663 665 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11514 662 670 663 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11513 7451 662 1168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11512 1168 662 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11511 3668 3743 3616 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11510 3616 3667 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11509 7451 3836 3668 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11508 3666 3668 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11507 7451 7095 7093 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11506 7092 7094 7091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11505 7091 7095 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11504 7091 7093 7092 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11503 7451 7090 7091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11502 7090 7094 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11501 7451 4368 2719 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11500 2719 2733 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11499 2719 4367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11498 7451 4724 2719 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11497 2718 2719 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11496 7451 4158 3924 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11495 3924 4161 4441 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11494 6992 6491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11493 5435 5833 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11492 3127 5377 3167 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11491 3126 5541 3127 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11490 7451 5378 3126 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11489 7451 6819 6679 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11488 6678 6676 6680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11487 6680 6819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11486 6680 6679 6678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11485 7451 6677 6680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11484 6677 6676 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11483 7451 3820 1840 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11482 1840 4934 4377 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11481 4985 5842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11480 7451 7108 4985 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11479 373 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11478 640 372 373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11477 371 953 640 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11476 7451 370 371 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_11475 4217 3636 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11474 7451 3637 4217 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11473 5954 5952 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11472 7451 5953 5954 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11471 5136 5369 5118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11470 5118 5134 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11469 7451 5226 5136 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11468 5282 5136 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11467 2692 3649 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11466 7451 2934 2691 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11465 7451 5128 2717 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11464 2716 5128 2692 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11463 2691 2717 2716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11462 2938 2716 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11461 5076 5074 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11460 7451 5075 5076 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11459 5600 5076 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11458 1106 5619 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11457 1106 4597 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11456 7451 1211 1106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11455 7451 1709 1106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11454 5885 3083 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11453 7451 3084 5885 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11452 5109 5127 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11451 7451 5125 5108 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11450 7451 5128 5131 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11449 5129 5128 5109 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11448 5108 5131 5129 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11447 5124 5129 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11446 3435 3804 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11445 7451 3475 3434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11444 7451 5128 3480 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11443 3479 5128 3435 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11442 3434 3480 3479 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11441 3476 3479 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11440 3437 4211 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11439 7451 3879 3436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11438 7451 5128 3493 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11437 3492 5128 3437 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11436 3436 3493 3492 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11435 3884 3492 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11434 3278 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11433 3321 4669 3278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11432 7451 3644 3321 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11431 2037 2814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11430 7451 2103 2037 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11429 1330 1334 1314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11428 1314 1333 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11427 7451 1332 1330 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11426 1552 1330 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11425 3738 3029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11424 3738 3037 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11423 7451 3033 3738 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11422 7451 3030 3738 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11421 4954 4996 4997 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11420 4955 5376 4954 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11419 4953 5087 4955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11418 7451 4995 4953 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11417 5819 4997 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11416 7451 7164 5117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11415 5117 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11414 5214 5137 5117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11413 5116 5275 5214 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11412 5117 5273 5116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11411 5620 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11410 5620 4441 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11409 7451 4448 5620 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11408 7451 4934 5620 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11407 1691 2926 1693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11406 1693 3135 1692 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11405 1692 3012 1693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11404 1691 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11403 7451 4979 1691 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11402 1693 6173 1691 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11401 1876 1692 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11400 7451 771 183 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11399 276 378 185 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11398 185 771 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11397 185 183 276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11396 7451 184 185 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11395 184 378 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11394 5265 5329 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11393 5331 6058 5265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11392 7451 5626 5331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11391 7451 6133 4085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11390 4085 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11389 4085 4158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11388 7451 7114 4085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11387 4084 4085 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11386 7451 1430 1350 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11385 1350 1723 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11384 1350 1466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11383 7451 2995 1350 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11382 2587 1350 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11381 7451 7164 5259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11380 5259 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11379 5411 5274 5259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11378 5258 5275 5411 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11377 5259 5273 5258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11376 498 609 538 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11375 496 495 498 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11374 497 847 496 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11373 7451 494 497 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11372 1841 538 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11371 5122 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11370 5299 5273 5122 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11369 7451 5887 5299 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11368 6140 6168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11367 6242 6169 6140 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11366 7451 6315 6242 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11365 6721 6751 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11364 6719 6752 6745 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11363 7451 7489 6719 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11362 6752 6753 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11361 7451 7215 6753 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11360 7451 6750 6751 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11359 6749 6752 6721 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11358 6720 6753 6749 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11357 7451 6746 6720 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11356 6746 6749 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11355 6745 6753 6746 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11354 7451 6745 7489 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11353 7489 6745 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11352 7451 2880 2268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11351 2268 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11350 7451 2881 2268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11349 2687 2268 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11348 6527 6560 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11347 6525 6556 6555 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11346 7451 7466 6525 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11345 6556 6557 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11344 7451 6528 6557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11343 7451 6561 6560 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11342 6559 6556 6527 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11341 6526 6557 6559 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11340 7451 6558 6526 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11339 6558 6559 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11338 6555 6557 6558 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11337 7451 6555 7466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11336 7466 6555 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11335 4765 4846 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11334 7451 4764 4765 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11333 4430 4986 4391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11332 4391 4581 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11331 7451 4427 4391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11330 4720 4430 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11329 4390 4987 4430 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11328 4391 4984 4390 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11327 4920 5137 4650 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11326 4650 5832 4920 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11325 7451 4649 4650 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11324 6144 6600 6179 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11323 6143 6599 6144 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11322 7451 6406 6143 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11321 6180 6179 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11320 5417 5418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11319 7451 6096 5417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11318 814 937 798 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11317 798 1728 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11316 7451 1681 814 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11315 1333 814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11314 5210 5207 5237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11313 5208 5818 5210 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11312 5209 5819 5208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11311 7451 5815 5209 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11310 5238 5237 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11309 4574 3411 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11308 7451 3412 4574 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11307 5227 5369 5228 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11306 5228 5225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11305 7451 5226 5227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11304 5806 5227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11303 4690 4718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11302 4722 5381 4690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11301 7451 6386 4722 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11300 2794 2847 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11299 7451 2846 2794 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11298 2748 1906 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11297 2748 1908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11296 7451 1915 2748 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11295 7451 2686 2748 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11294 6568 7042 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11293 6568 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11292 7451 5746 6568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11291 7451 7114 6568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11290 3217 3216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11289 7451 6894 3217 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11288 3304 3217 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11287 550 4161 1051 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11286 606 4934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11285 7451 606 550 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11284 7203 7379 7204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11283 7204 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11282 7451 7475 7203 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11281 7419 7203 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11280 7451 1355 1321 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11279 1321 1356 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11278 1872 2502 1321 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11277 1320 2435 1872 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11276 1321 2853 1320 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11275 1329 1444 1383 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11274 1328 1508 1329 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11273 7451 1627 1328 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_11272 1382 1383 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11271 4373 6600 4372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11270 4371 4514 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11269 7451 4371 4373 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11268 7451 3633 2998 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11267 2998 2999 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11266 2998 3632 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11265 7451 3300 2998 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11264 3216 2998 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11263 5382 5457 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11262 7451 6333 5382 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11261 6979 5382 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11260 7451 2222 2223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11259 2223 2418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11258 7451 2220 2223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11257 2221 2223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11256 2442 2664 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11255 3005 5882 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11254 7451 1558 1349 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11253 1550 1427 1319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11252 1319 1558 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11251 1319 1349 1550 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11250 7451 1347 1319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11249 1347 1427 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11248 7451 4437 3999 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11247 3999 4081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11246 3999 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11245 7451 7162 3999 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11244 4511 3999 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11243 7451 2111 813 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11242 813 2602 5173 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11241 5207 5160 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11240 2517 2934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11239 4838 5137 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11238 2127 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11237 2165 2929 2127 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11236 7451 5882 2165 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11235 3748 3783 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11234 3746 3782 3776 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11233 7451 3774 3746 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11232 3782 3784 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11231 7451 4638 3784 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11230 7451 3779 3783 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11229 3780 3782 3748 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11228 3747 3784 3780 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11227 7451 3777 3747 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11226 3777 3780 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11225 3776 3784 3777 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11224 7451 3776 3774 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11223 3774 3776 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11222 2825 2688 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11221 7451 2687 2825 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11220 4628 4752 4629 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11219 4627 4833 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11218 7451 4627 4628 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11217 7451 7418 7415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11216 7416 7465 7417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11215 7417 7418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11214 7417 7415 7416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11213 7451 7414 7417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11212 7414 7465 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11211 1287 1577 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11210 7451 5000 1287 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11209 5723 5505 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11208 7451 5506 5723 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11207 3084 2659 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11206 7451 2707 3084 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11205 2806 3649 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11204 7451 3086 2804 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11203 7451 4106 2807 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11202 2805 4106 2806 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11201 2804 2807 2805 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11200 3092 2805 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11199 4087 5127 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11198 7451 4104 4086 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11197 7451 4106 4109 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11196 4108 4106 4087 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11195 4086 4109 4108 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11194 4103 4108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11193 1896 2814 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11192 7451 2811 1896 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11191 3699 3804 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11190 7451 3696 3697 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11189 7451 4106 3700 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11188 3698 4106 3699 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11187 3697 3700 3698 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11186 3695 3698 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11185 3707 4211 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11184 7451 4113 3706 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11183 7451 4106 3709 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11182 3708 4106 3707 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11181 3706 3709 3708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11180 4119 3708 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11179 4922 4920 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11178 7451 4921 4922 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11177 5521 4922 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11176 6399 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11175 6399 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11174 7451 5969 6399 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11173 7451 7114 6399 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11172 7451 7390 5544 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11171 7451 7388 5545 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11170 5544 5545 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11169 7451 5994 2824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11168 2824 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11167 2823 6266 2824 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11166 2822 5840 2823 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11165 2824 6332 2822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11164 7123 7431 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11163 7451 7107 7123 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11162 834 832 807 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11161 807 960 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11160 7451 2592 834 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11159 833 834 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11158 1260 1547 1259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11157 1259 1732 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11156 7451 1548 1260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11155 2007 1260 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11154 3124 3129 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11153 3131 4695 3124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11152 7451 3128 3131 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11151 6007 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11150 6042 6566 6007 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11149 7451 6676 6042 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11148 6429 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11147 6471 7228 6429 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11146 7451 7466 6471 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11145 7451 6843 6132 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11144 6132 6405 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11143 6132 6768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11142 7451 6907 6132 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11141 7034 6132 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11140 6095 6372 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11139 6094 6293 6095 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11138 7451 7420 6094 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11137 6146 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11136 6185 7228 6146 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11135 7451 7493 6185 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11134 7451 7074 6867 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11133 7011 7453 6856 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11132 6856 7074 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11131 6856 6867 7011 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11130 7451 6865 6856 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11129 6865 7453 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11128 6 39 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11127 4 38 33 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11126 7451 6266 4 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11125 38 40 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11124 7451 403 40 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11123 7451 41 39 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11122 36 38 6 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11121 5 40 36 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11120 7451 34 5 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11119 34 36 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11118 33 40 34 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11117 7451 33 6266 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11116 6266 33 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11115 5094 5844 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11114 7451 5889 5094 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11113 5093 5094 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11112 2186 2183 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11111 7451 2182 2186 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11110 2185 2186 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11109 1904 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11108 7451 1976 1904 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11107 2322 1904 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11106 7451 3890 3765 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11105 3765 4228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11104 7105 3814 3765 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11103 3764 4149 7105 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11102 3765 5909 3764 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11101 2277 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11100 2508 2929 2277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11099 7451 6025 2508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11098 7451 2514 2096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11097 2096 2383 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11096 7451 2304 2096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11095 2095 2096 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11094 7451 4156 4157 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11093 7451 4158 4160 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11092 4157 4160 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11091 5911 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11090 7451 7384 5911 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11089 5909 5911 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11088 6717 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11087 6731 7428 6717 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11086 7451 6965 6731 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11085 929 972 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11084 927 971 964 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11083 7451 963 927 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11082 971 973 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11081 7451 1290 973 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11080 7451 968 972 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11079 969 971 929 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11078 928 973 969 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11077 7451 966 928 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11076 966 969 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11075 964 973 966 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11074 7451 964 963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11073 963 964 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11072 3426 3742 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11071 3732 3425 3426 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11070 7451 4148 3732 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11069 6139 6166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11068 6593 6165 6139 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11067 7451 6315 6593 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11066 7451 4568 1969 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11065 1969 2452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11064 1969 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11063 7451 4569 1969 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11062 1968 1969 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11061 7451 4161 2399 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11060 2399 2602 2684 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11059 1167 2541 1166 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11058 1166 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11057 7451 1445 1167 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11056 1837 1167 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11055 4175 4305 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11054 7451 4175 4173 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_11053 4174 4172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11052 7451 4174 4102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11051 4102 4173 4170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11050 4170 4175 4101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11049 4100 4937 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11048 7451 4166 4937 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11047 4937 4166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11046 4101 4167 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11045 4167 4170 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11044 7451 7500 4167 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11043 4166 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_11042 4166 4173 4100 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11041 4167 4175 4166 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_11040 4774 5072 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11039 7451 4773 4774 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11038 6843 7114 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11037 6843 5994 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11036 7451 6133 6843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11035 7451 6981 6583 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11034 6584 6599 6968 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11033 6585 6848 6584 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11032 6583 6600 6585 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_11031 4970 5369 4942 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11030 4942 4971 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11029 7451 5226 4970 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11028 5801 4970 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11027 2658 3213 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11026 7451 2657 2658 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11025 1442 1440 1443 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11024 1443 1441 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11023 7451 4597 1442 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11022 1759 1442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11021 844 1908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11020 7451 1915 844 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11019 7451 2686 3425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11018 7451 4934 2611 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11017 3425 2611 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_11016 3812 4360 3763 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11015 3763 3811 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11014 7451 6041 3812 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11013 3810 3812 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11012 6023 7462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11011 6023 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11010 7451 6968 6023 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11009 7152 7428 7121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11008 7121 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11007 7451 7493 7152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11006 7151 7152 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_11005 2608 7162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11004 2608 2390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11003 7451 2255 2608 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11002 4230 4297 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11001 7451 4588 4230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_11000 4231 4230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10999 1063 2842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10998 1082 2792 1063 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10997 7451 2133 1082 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10996 2155 2434 2126 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10995 2126 2154 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10994 7451 2164 2155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10993 2153 2155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10992 4588 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10991 4588 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10990 7451 4437 4588 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10989 7451 7114 4588 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10988 6839 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10987 6839 6914 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10986 7451 7164 6839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10985 7451 7113 6839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10984 7451 5079 5080 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10983 5080 6832 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10982 7451 5238 5080 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10981 5078 5080 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10980 1767 1906 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10979 1767 1908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10978 7451 1915 1767 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10977 7451 4000 1767 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10976 4569 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10975 4569 1292 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10974 7451 4081 4569 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10973 7451 5690 4569 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10972 5997 6061 7384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10971 5996 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10970 7451 5996 5997 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10969 2085 2524 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10968 2085 2141 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10967 7451 4694 2085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10966 7451 2228 2085 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10965 7451 6193 6050 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10964 6050 6048 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10963 7451 6046 6050 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10962 6047 6050 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10961 7451 7164 7167 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10960 7167 7391 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10959 7451 7162 7167 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10958 7163 7167 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10957 6093 6118 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10956 6091 6120 6115 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10955 7451 7452 6091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10954 6120 6121 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10953 7451 6231 6121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10952 7451 6119 6118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10951 6117 6120 6093 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10950 6092 6121 6117 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10949 7451 6116 6092 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10948 6116 6117 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10947 6115 6121 6116 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10946 7451 6115 7452 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10945 7452 6115 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10944 4503 4502 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10943 4649 5381 4503 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10942 7451 6386 4649 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10941 2703 4695 2689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10940 2689 3149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10939 7451 3213 2703 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10938 2847 2703 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10937 7451 3167 472 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10936 434 472 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10935 7451 472 434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10934 7451 472 434 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10933 434 472 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10932 7451 434 386 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10931 1688 386 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10930 7451 386 1688 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10929 7451 386 1688 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10928 1688 386 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10927 7451 434 328 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10926 3546 328 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10925 7451 328 3546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10924 7451 328 3546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10923 3546 328 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10922 7451 579 285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10921 331 285 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10920 7451 285 331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10919 7451 285 331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10918 331 285 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10917 7451 331 332 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10916 3352 332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10915 7451 332 3352 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10914 7451 332 3352 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10913 3352 332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10912 7451 331 228 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10911 4934 228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10910 7451 228 4934 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10909 7451 228 4934 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10908 4934 228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10907 5853 5872 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10906 5851 5875 5866 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10905 7451 6628 5851 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10904 5875 5874 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10903 7451 6302 5874 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10902 7451 5870 5872 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10901 5871 5875 5853 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10900 5852 5874 5871 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10899 7451 5868 5852 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10898 5868 5871 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10897 5866 5874 5868 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10896 7451 5866 6628 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10895 6628 5866 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10894 2283 3837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10893 2456 2467 2283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10892 2282 2338 2456 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10891 7451 2337 2282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_10890 6517 6543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10889 6515 6544 6540 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10888 7451 6539 6515 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10887 6544 6545 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10886 7451 6622 6545 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10885 7451 6549 6543 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10884 6542 6544 6517 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10883 6516 6545 6542 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10882 7451 6546 6516 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10881 6546 6542 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10880 6540 6545 6546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10879 7451 6540 6539 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10878 6539 6540 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10877 2128 3214 4697 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10876 2167 2168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10875 7451 2167 2128 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10874 4696 4104 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10873 5134 4834 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10872 3771 6432 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10871 6536 6714 6538 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10870 6537 6852 6536 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10869 7451 7113 6537 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10868 1198 1823 1174 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10867 1174 1287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10866 7451 1197 1198 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10865 2029 1198 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10864 2402 2449 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10863 2400 2450 2444 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10862 7451 2602 2400 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10861 2450 2451 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10860 7451 2533 2451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10859 7451 2603 2449 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10858 2446 2450 2402 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10857 2401 2451 2446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10856 7451 2445 2401 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10855 2445 2446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10854 2444 2451 2445 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10853 7451 2444 2602 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10852 2602 2444 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10851 5653 5969 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10850 4112 6175 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10849 7451 5171 5170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10848 5170 5172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10847 5170 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10846 7451 6266 5170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10845 5457 5170 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10844 3874 4908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10843 3877 4413 3874 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10842 3873 4411 3877 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10841 7451 4197 3873 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10840 3878 3877 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10839 7451 3352 912 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10838 912 4158 2392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10837 495 4517 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10836 7451 405 495 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10835 7451 3979 1712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10834 1712 1727 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10833 1728 3546 1712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10832 1711 2139 1728 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10831 1712 1866 1711 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10830 5960 5809 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10829 7451 5877 5960 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10828 7079 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10827 7078 7428 7079 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10826 7451 7453 7078 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10825 3386 3387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10824 7451 4504 3385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10823 7451 4264 3388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10822 3417 4264 3386 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10821 3385 3388 3417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10820 3582 3417 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10819 5127 3470 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10818 5127 3472 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10817 7451 3469 5127 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10816 3122 3410 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10815 7451 4502 3121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10814 7451 4264 3153 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10813 3151 4264 3122 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10812 3121 3153 3151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10811 3315 3151 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10810 4241 4265 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10809 7451 4716 4242 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10808 7451 4264 4267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10807 4263 4264 4241 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10806 4242 4267 4263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10805 4261 4263 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10804 951 1435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10803 951 1968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10802 7451 1700 951 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10801 4829 4828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10800 7451 6266 4829 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10799 2416 2508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10798 2416 3769 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10797 7451 2507 2416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10796 2877 4372 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10795 7451 3347 2877 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10794 2875 2877 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10793 3439 3495 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10792 7451 4861 3438 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10791 7451 4264 3498 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10790 3497 4264 3439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10789 3438 3498 3497 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10788 3797 3497 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10787 1815 3546 1816 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10786 1816 1869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10785 7451 3000 1816 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10784 1813 1815 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10783 1814 2095 1815 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10782 1816 1866 1814 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10781 3744 4446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10780 3744 5172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10779 7451 5173 3744 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10778 7451 3742 3744 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10777 7451 6094 5661 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10776 5661 5660 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10775 7451 5803 5661 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10774 5659 5661 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10773 2947 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10772 2948 2946 2947 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10771 7451 5055 2948 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10770 6572 7042 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10769 6572 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10768 7451 6187 6572 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10767 7451 6333 6572 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10766 1045 1837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10765 7451 7114 1045 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10764 1044 1045 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10763 5986 5985 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10762 7451 6181 5986 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10761 5984 5986 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10760 1964 6173 1963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10759 2159 3012 1964 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10758 1964 3135 2159 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10757 1963 2926 1964 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10756 1963 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10755 7451 4979 1963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10754 7451 5835 5836 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10753 5836 6328 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10752 7451 6471 5836 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10751 5834 5836 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10750 1189 2792 1173 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10749 1173 2842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10748 7451 2133 1189 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10747 1187 1189 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10746 1706 1833 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10745 7451 7114 1706 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10744 2035 1706 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10743 7451 6979 6842 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10742 6842 6980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10741 7451 7480 6842 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10740 6841 6842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10739 7451 6705 6706 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10738 6706 6764 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10737 7451 6899 6706 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10736 6704 6706 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10735 5257 6166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10734 5503 6165 5257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10733 7451 5876 5503 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10732 6692 6691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10731 6686 6695 6685 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10730 7451 7494 6686 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10729 6695 6694 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10728 7451 6693 6694 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10727 7451 6690 6691 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10726 6688 6695 6692 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10725 6689 6694 6688 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10724 7451 6687 6689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10723 6687 6688 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10722 6685 6694 6687 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10721 7451 6685 7494 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10720 7494 6685 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10719 7451 7477 7368 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10718 7372 7369 7346 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10717 7346 7477 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10716 7346 7368 7372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10715 7451 7371 7346 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10714 7371 7369 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10713 5697 6168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10712 5738 6169 5697 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10711 7451 5815 5738 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10710 7451 5171 1165 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10709 1165 1775 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10708 7451 2881 1165 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10707 1501 1165 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10706 4791 5691 4792 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10705 4792 5842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10704 7451 6133 4791 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10703 4790 4791 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10702 2830 2846 2831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10701 2831 2991 2849 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10700 2849 2995 2831 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10699 2830 2931 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10698 7451 4254 2830 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10697 2831 2847 2830 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10696 2844 2849 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10695 7451 1149 1027 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10694 1146 1732 1028 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10693 1028 1149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10692 1028 1027 1146 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10691 7451 1026 1028 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10690 1026 1732 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10689 6953 6975 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10688 6951 6977 6971 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10687 7451 7480 6951 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10686 6977 6974 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10685 7451 7225 6974 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10684 7451 6976 6975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10683 6973 6977 6953 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10682 6952 6974 6973 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10681 7451 6972 6952 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10680 6972 6973 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10679 6971 6974 6972 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10678 7451 6971 7480 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10677 7480 6971 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10676 5229 5230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10675 7451 5366 5229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10674 2810 3810 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10673 7451 3013 2810 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10672 3119 5000 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10671 3119 5994 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10670 7451 6133 3119 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10669 571 3546 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10668 571 771 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10667 7451 1082 571 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10666 2102 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10665 2102 1570 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10664 7451 2033 2102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10663 7451 5690 2102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10662 6599 6046 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10661 6599 6193 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10660 7451 6048 6599 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10659 4773 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10658 4773 4081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10657 7451 4437 4773 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10656 7451 7162 4773 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10655 7451 280 220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10654 372 276 200 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10653 200 280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10652 200 220 372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10651 7451 218 200 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10650 218 276 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10649 7451 6162 5808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10648 5808 5806 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10647 7451 5807 5808 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10646 5805 5808 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10645 1717 1750 1716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10644 2865 1880 1717 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10643 1717 1876 2865 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10642 1716 1749 1717 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10641 1716 1746 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10640 7451 1747 1716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10639 6834 6886 6835 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10638 6835 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10637 7451 7034 6835 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10636 6832 6834 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10635 6833 7032 6834 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10634 6835 7313 6833 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10633 7451 6332 5689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10632 5689 6266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10631 7451 7114 5689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10630 5688 5689 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10629 5309 5306 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10628 7451 5897 5309 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10627 5307 5309 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10626 3414 3636 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10625 7451 3637 3414 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10624 3495 3414 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10623 3408 3407 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10622 7451 3406 3408 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10621 3562 3408 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10620 1160 2816 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10619 7451 1577 1160 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10618 1159 1160 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10617 5070 5735 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10616 5421 5734 5070 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10615 7451 5069 5421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10614 4287 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10613 7451 4589 4287 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10612 4583 4287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10611 1088 1768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10610 7451 1435 1088 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10609 1466 1088 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10608 551 3546 540 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10607 540 2290 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10606 7451 3625 540 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10605 1636 551 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10604 539 3549 551 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10603 540 1866 539 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10602 3234 4066 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10601 7451 3322 3234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10600 3233 3234 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10599 6844 7109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10598 7451 7042 6844 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10597 7334 6844 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10596 986 5171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10595 7451 1775 986 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10594 4437 986 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10593 2143 2292 2124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10592 2124 3023 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10591 7451 2392 2124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10590 2140 2143 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10589 2123 2141 2143 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10588 2124 2139 2123 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10587 7451 1968 954 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10586 954 2718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10585 954 1700 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10584 7451 1688 954 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10583 953 954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10582 4971 5274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10581 3129 3868 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10580 3149 3774 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10579 4841 5055 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10578 3481 3696 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10577 7451 4081 111 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10576 111 4437 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10575 7451 6266 111 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10574 195 111 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10573 7451 1548 1172 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10572 1172 1952 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10571 1182 1337 1172 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10570 1171 1419 1182 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10569 1172 1336 1171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10568 7451 4377 4374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10567 4374 4447 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10566 4374 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10565 7451 4376 4374 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10564 7109 4374 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10563 2274 2288 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10562 3070 2287 2274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10561 7451 2784 3070 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10560 6613 6614 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10559 7451 6851 6613 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10558 5913 5912 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10557 7451 7162 5913 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10556 5504 6316 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10555 5953 6314 5504 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10554 7451 5876 5953 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10553 6648 7496 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10552 6648 7164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10551 7451 7286 6648 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10550 5368 5884 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10549 5675 5885 5368 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10548 7451 5815 5675 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10547 7451 1034 1035 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10546 5884 1032 1033 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10545 1033 1034 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10544 1033 1035 5884 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10543 7451 1031 1033 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10542 1031 1032 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10541 2982 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10540 3013 4669 2982 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10539 7451 3012 3013 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10538 2926 4569 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10537 2926 4568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10536 7451 4588 2926 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10535 935 2111 1915 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10534 988 2602 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10533 7451 988 935 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10532 6409 6407 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10531 6409 6710 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10530 7451 6906 6409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10529 7451 6408 6409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10528 3282 4987 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10527 3649 4984 3282 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10526 7451 4986 3649 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10525 7142 7428 7118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10524 7118 7280 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10523 7451 7466 7142 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10522 7210 7142 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10521 3585 3581 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10520 7451 3585 3583 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10519 3584 3582 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10518 7451 3584 3580 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10517 3580 3583 3579 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10516 3579 3585 3578 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10515 3575 4504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10514 7451 3576 4504 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10513 4504 3576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10512 3578 3577 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10511 3577 3579 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10510 7451 7500 3577 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10509 3576 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10508 3576 3583 3575 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10507 3577 3585 3576 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10506 5074 5216 4770 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10505 4770 5832 5074 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10504 7451 4769 4770 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10503 1491 1489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10502 7451 1694 1491 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10501 3160 1491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10500 6331 7164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10499 7451 7286 6331 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10498 6981 6331 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10497 4666 4995 4780 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10496 4665 4726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10495 7451 4665 4666 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10494 4369 4368 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10493 7451 4367 4369 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10492 4781 4369 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10491 3421 4568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10490 7451 4569 3421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10489 3420 3421 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10488 6281 6757 6326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10487 6324 6325 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10486 7451 6324 6281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10485 1157 2435 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10484 1197 2853 1157 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10483 7451 2504 1197 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10482 7451 6332 6265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10481 6265 7042 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10480 7451 7162 6265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10479 6338 6265 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10478 2941 2942 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10477 2935 2943 2936 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10476 7451 2934 2935 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10475 2943 2944 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10474 7451 3571 2944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10473 7451 2938 2942 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10472 2940 2943 2941 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10471 2939 2944 2940 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10470 7451 2937 2939 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10469 2937 2940 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10468 2936 2944 2937 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10467 7451 2936 2934 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10466 2934 2936 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10465 5107 5554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10464 7451 5107 5106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10463 5105 5393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10462 7451 5105 5104 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10461 5104 5106 5103 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10460 5103 5107 5102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10459 5098 7388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10458 7451 5099 7388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10457 7388 5099 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10456 5102 5101 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10455 5101 5103 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10454 7451 5100 5101 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10453 5099 5100 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10452 5099 5106 5098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10451 5101 5107 5099 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10450 4907 6316 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10449 5352 6314 4907 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10448 7451 5069 5352 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10447 5974 5711 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10446 7451 5738 5974 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10445 7451 6061 5845 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10444 5845 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10443 5845 7390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10442 7451 7388 5845 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10441 5912 5845 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10440 1315 1333 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10439 1420 1334 1315 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10438 7451 1332 1420 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10437 7451 2082 2005 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10436 5735 2002 1983 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10435 1983 2082 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10434 1983 2005 5735 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10433 7451 2003 1983 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10432 2003 2002 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10431 3430 3922 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10430 3736 3925 3430 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10429 7451 5055 3736 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10428 2180 2541 2129 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10427 2129 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10426 7451 2179 2180 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10425 2390 2180 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10424 2219 2221 3472 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10423 2218 2366 2219 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10422 7451 2217 2218 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10421 6956 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10420 6955 7228 6956 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10419 7451 7464 6955 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10418 4857 5078 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10417 7451 4720 4857 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10416 6202 6135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10415 6202 6410 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10414 7451 6992 6202 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10413 5965 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10412 6124 7379 5965 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10411 7451 6676 6124 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10410 6141 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10409 6306 6394 6141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10408 7451 6173 6306 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10407 6837 7480 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10406 6837 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10405 7451 6968 6837 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10404 2854 3135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10403 7451 3645 2854 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10402 5407 5467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10401 5468 5466 5407 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10400 5406 5695 5468 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10399 7451 5544 5406 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10398 6056 5468 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10397 446 1304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10396 446 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10395 7451 3346 446 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10394 239 1906 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10393 239 2887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10392 7451 3346 239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10391 5985 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10390 5985 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10389 7451 5536 5985 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10388 7451 7162 5985 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10387 2710 4695 2690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10386 2690 3710 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10385 7451 3145 2710 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10384 2800 2710 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_10383 7451 3655 3656 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10382 4074 5138 3619 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10381 3619 3655 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10380 3619 3656 4074 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10379 7451 3653 3619 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10378 3653 5138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10377 7451 7489 7096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10376 7096 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10375 7451 7494 7096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10374 7095 7096 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10373 5814 6166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10372 5813 6165 5814 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10371 7451 5815 5813 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10370 2409 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10369 2521 2946 2409 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10368 7451 4834 2521 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10367 801 1146 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10366 1547 1182 801 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10365 7451 1145 1547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10364 6381 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10363 6380 7379 6381 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10362 7451 6628 6380 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10361 5658 5724 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10360 5656 5725 5721 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10359 7451 7454 5656 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10358 5725 5726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10357 7451 6231 5726 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10356 7451 5723 5724 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10355 5706 5725 5658 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10354 5657 5726 5706 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10353 7451 5705 5657 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10352 5705 5706 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10351 5721 5726 5705 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10350 7451 5721 7454 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10349 7454 5721 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10348 947 949 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10347 7451 951 947 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10346 1145 947 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10345 6129 6128 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10344 7451 6402 6129 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10343 6325 6129 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10342 7451 1914 1850 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10341 1850 1911 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10340 2325 2536 1850 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10339 1849 2398 2325 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10338 1850 2813 1849 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10337 2251 4161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10336 7451 2602 2251 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10335 2811 2251 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10334 6995 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10333 7016 7379 6995 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10332 7451 7462 7016 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10331 5796 5798 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10330 5791 5799 5792 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10329 7451 6965 5791 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10328 5799 5800 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10327 7451 6231 5800 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10326 7451 5797 5798 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10325 5794 5799 5796 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10324 5795 5800 5794 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10323 7451 5793 5795 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10322 5793 5794 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10321 5792 5800 5793 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10320 7451 5792 6965 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10319 6965 5792 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10318 7451 1968 1226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10317 1226 1700 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10316 7451 1435 1226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10315 1866 1226 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10314 7451 6726 6228 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10313 6226 7335 6227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10312 6227 6726 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10311 6227 6228 6226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10310 7451 6225 6227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10309 6225 7335 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10308 4941 4968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10307 4939 4967 4961 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10306 7451 4959 4939 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10305 4967 4969 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10304 7451 5584 4969 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10303 7451 4966 4968 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10302 4963 4967 4941 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10301 4940 4969 4963 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10300 7451 4962 4940 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10299 4962 4963 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10298 4961 4969 4962 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10297 7451 4961 4959 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10296 4959 4961 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10295 7451 4207 4099 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10294 4099 4228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10293 5989 4148 4099 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10292 4098 4149 5989 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10291 4099 5909 4098 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10290 7451 1304 1050 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10289 1050 1906 1440 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10288 7465 7464 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10287 4412 6035 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10286 5371 5536 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10285 7451 3210 3133 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10284 3132 3133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10283 7451 3133 3132 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10282 7451 3133 3132 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10281 3132 3133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10280 7451 3210 3205 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10279 3204 3205 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10278 7451 3205 3204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10277 7451 3205 3204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10276 3204 3205 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10275 7451 3210 3206 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10274 3400 3206 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10273 7451 3206 3400 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10272 7451 3206 3400 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10271 3400 3206 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10270 7451 3210 3141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10269 3140 3141 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10268 7451 3141 3140 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10267 7451 3141 3140 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10266 3140 3141 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10265 7451 3210 3209 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10264 3208 3209 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10263 7451 3209 3208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10262 7451 3209 3208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10261 3208 3209 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10260 7451 3210 3211 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10259 3558 3211 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10258 7451 3211 3558 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10257 7451 3211 3558 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10256 3558 3211 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10255 7451 3229 2152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10254 2151 2152 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10253 7451 2152 2151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10252 7451 2152 2151 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10251 2151 2152 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10250 2693 2926 2694 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10249 2694 3135 2700 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10248 2700 3644 2694 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10247 2693 2925 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10246 7451 5216 2693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10245 2694 6388 2693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10244 2696 2700 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10243 6733 6676 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10242 3811 3727 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10241 5837 5616 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10240 7451 5457 5837 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10239 6561 6309 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10238 7451 6246 6561 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10237 7451 3229 2233 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10236 2232 2233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10235 7451 2233 2232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10234 7451 2233 2232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10233 2232 2233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10232 7451 3229 2235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10231 2234 2235 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10230 7451 2235 2234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10229 7451 2235 2234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10228 2234 2235 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10227 7451 3229 2162 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10226 2163 2162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10225 7451 2162 2163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10224 7451 2162 2163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10223 2163 2162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10222 7451 3229 2238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10221 2237 2238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10220 7451 2238 2237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10219 7451 2238 2237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10218 2237 2238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10217 7451 3229 2240 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10216 2239 2240 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10215 7451 2240 2239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10214 7451 2240 2239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10213 2239 2240 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10212 7451 3229 3148 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10211 3147 3148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10210 7451 3148 3147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10209 7451 3148 3147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10208 3147 3148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10207 7451 3229 3219 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10206 3218 3219 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10205 7451 3219 3218 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10204 7451 3219 3218 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10203 3218 3219 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10202 7451 3229 3221 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10201 3220 3221 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10200 7451 3221 3220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10199 7451 3221 3220 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10198 3220 3221 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10197 7451 7477 7277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10196 7274 7480 7250 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10195 7250 7477 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10194 7250 7277 7274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10193 7451 7273 7250 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10192 7273 7480 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10191 2505 2785 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10190 7451 2837 2505 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10189 7451 6852 6716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10188 6716 6714 6715 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10187 6849 6715 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10186 5822 5817 5823 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10185 5820 5818 5822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10184 5821 5819 5820 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10183 7451 5815 5821 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_10182 5816 5823 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10181 7451 5600 5601 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10180 5601 6637 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10179 7451 5669 5601 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10178 5711 5601 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10177 3266 5691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10176 7451 5001 3266 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10175 2653 2507 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10174 2653 2583 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10173 7451 3769 2653 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10172 7451 2508 2653 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10171 7451 3229 3154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10170 3155 3154 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10169 7451 3154 3155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10168 7451 3154 3155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10167 3155 3154 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10166 7451 3229 3228 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10165 3227 3228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10164 7451 3228 3227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10163 7451 3228 3227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10162 3227 3228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10161 7451 3229 3230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10160 3571 3230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10159 7451 3230 3571 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10158 7451 3230 3571 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10157 3571 3230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10156 7451 2712 852 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10155 1264 852 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10154 7451 852 1264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10153 7451 852 1264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10152 1264 852 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10151 1835 1906 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10150 1835 1908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10149 7451 1915 1835 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10148 1055 3820 4448 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10147 1054 4376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10146 7451 1054 1055 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10145 7451 7235 6344 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10144 7451 6652 5995 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10143 6344 5995 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_10142 1216 1543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10141 1216 266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10140 7451 1025 1216 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10139 1689 1688 1690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10138 1690 1876 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10137 7451 1851 1690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10136 1686 1689 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10135 1687 2095 1689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10134 1690 3545 1687 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10133 7451 7335 6870 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10132 6870 7074 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10131 6870 7452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10130 7451 7453 6870 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10129 6869 6870 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10128 7451 2712 856 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10127 1281 856 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10126 7451 856 1281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10125 7451 856 1281 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10124 1281 856 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10123 7451 2712 2701 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10122 3210 2701 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10121 7451 2701 3210 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10120 7451 2701 3210 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10119 3210 2701 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10118 7451 2712 2713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10117 3229 2713 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10116 7451 2713 3229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10115 7451 2713 3229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10114 3229 2713 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10113 7120 7151 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10112 7149 7315 7120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10111 7451 7420 7149 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10110 4053 4488 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10109 7451 4053 4054 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_10108 4052 4261 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10107 7451 4052 4051 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10106 4051 4054 4048 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10105 4048 4053 4049 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10104 4046 4716 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10103 7451 4047 4716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10102 4716 4047 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10101 4049 4050 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10100 4050 4048 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10099 7451 7500 4050 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10098 4047 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_10097 4047 4054 4046 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10096 4050 4053 4047 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_10095 3600 3922 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10094 3601 3925 3600 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10093 7451 5274 3601 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10092 7451 1295 330 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10091 329 330 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10090 7451 330 329 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10089 7451 330 329 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10088 329 330 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10087 7451 1295 388 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10086 387 388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10085 7451 388 387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10084 7451 388 387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10083 387 388 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10082 7451 1295 389 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10081 788 389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10080 7451 389 788 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10079 7451 389 788 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10078 788 389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10077 7451 1295 334 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10076 333 334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10075 7451 334 333 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10074 7451 334 333 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10073 333 334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10072 7451 1295 393 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10071 392 393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10070 7451 393 392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10069 7451 393 392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10068 392 393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10067 7451 1295 394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10066 598 394 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10065 7451 394 598 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10064 7451 394 598 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10063 598 394 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10062 7451 1295 1230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10061 1201 1230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10060 7451 1230 1201 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10059 7451 1230 1201 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10058 1201 1230 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10057 3721 4142 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10056 7451 3719 3721 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10055 3720 3721 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10054 1162 1365 1163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10053 1163 1368 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10052 7451 4437 1163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10051 1971 1162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10050 1161 1366 1162 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10049 1163 1500 1161 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10048 2389 4934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10047 7451 4158 2389 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10046 2816 2389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10045 7336 7390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10044 7451 7388 7336 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10043 7353 7336 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10042 917 1109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10041 7451 1111 917 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_10040 1620 917 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10039 3215 3214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10038 3213 3212 3215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10037 7451 3550 3213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10036 7451 1295 1289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10035 1288 1289 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10034 7451 1289 1288 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10033 7451 1289 1288 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10032 1288 1289 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10031 7451 1295 1291 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10030 1290 1291 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10029 7451 1291 1290 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10028 7451 1291 1290 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10027 1290 1291 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10026 7451 1295 1234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10025 1206 1234 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10024 7451 1234 1206 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10023 7451 1234 1206 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10022 1206 1234 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10021 7451 1295 1293 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10020 1294 1293 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10019 7451 1293 1294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10018 7451 1293 1294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10017 1294 1293 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10016 7451 1295 1297 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10015 1296 1297 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10014 7451 1297 1296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10013 7451 1297 1296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10012 1296 1297 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10011 7451 1310 336 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10010 335 336 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10009 7451 336 335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10008 7451 336 335 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10007 335 336 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10006 7451 1310 397 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10005 396 397 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10004 7451 397 396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10003 7451 397 396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10002 396 397 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10001 7451 1310 398 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_10000 669 398 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09999 7451 398 669 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09998 7451 398 669 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09997 669 398 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09996 4533 4560 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09995 4531 4562 4555 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09994 7451 6173 4531 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09993 4562 4563 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09992 7451 4561 4563 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09991 7451 4644 4560 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09990 4557 4562 4533 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09989 4532 4563 4557 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09988 7451 4556 4532 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09987 4556 4557 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09986 4555 4563 4556 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09985 7451 4555 6173 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09984 6173 4555 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09983 7451 4600 1042 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09982 1042 1292 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09981 1042 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09980 7451 5690 1042 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09979 1569 1042 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09978 7451 1581 1378 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09977 1378 1631 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09976 1378 1377 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09975 7451 1618 1378 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09974 1376 1378 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09973 7451 1292 532 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09972 532 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09971 7451 6266 532 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09970 533 532 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09969 2538 2541 2539 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09968 2539 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09967 7451 2542 2538 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09966 2537 2538 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09965 6850 7287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09964 6848 6849 6850 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09963 6847 6845 6848 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09962 7451 6846 6847 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09961 7451 5171 4936 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09960 4936 5172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09959 4936 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09958 7451 6133 4936 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09957 6565 4936 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09956 4606 5691 4540 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09955 4540 5842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09954 7451 5841 4606 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09953 4604 4606 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09952 6106 6314 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09951 7107 6316 6106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09950 7451 6125 7107 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09949 7451 1310 344 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09948 343 344 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09947 7451 344 343 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09946 7451 344 343 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09945 343 344 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09944 7451 1310 402 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09943 401 402 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09942 7451 402 401 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09941 7451 402 401 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09940 401 402 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09939 7451 1310 404 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09938 403 404 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09937 7451 404 403 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09936 7451 404 403 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09935 403 404 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09934 7451 1310 1238 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09933 1210 1238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09932 7451 1238 1210 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09931 7451 1238 1210 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09930 1210 1238 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09929 7451 1310 1301 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09928 1300 1301 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09927 7451 1301 1300 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09926 7451 1301 1300 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09925 1300 1301 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09924 7451 1310 1303 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09923 1302 1303 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09922 7451 1303 1302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09921 7451 1303 1302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09920 1302 1303 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09919 7451 1310 1244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09918 1215 1244 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09917 7451 1244 1215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09916 7451 1244 1215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09915 1215 1244 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09914 4689 4716 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09913 4769 5381 4689 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09912 7451 6386 4769 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09911 2168 1568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09910 7451 1569 2168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09909 4076 4589 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09908 5012 4074 4076 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09907 7451 4075 5012 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09906 4840 5369 4795 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09905 4795 4838 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09904 7451 5226 4840 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09903 5728 4840 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09902 7444 7508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09901 7451 7444 7443 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09900 7442 7440 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09899 7451 7442 7441 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09898 7441 7443 7439 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09897 7439 7444 7438 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09896 7435 7512 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09895 7451 7436 7512 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09894 7512 7436 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09893 7438 7437 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09892 7437 7439 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09891 7451 7500 7437 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09890 7436 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09889 7436 7443 7435 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09888 7437 7444 7436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_09887 5429 5520 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09886 7451 5813 5429 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09885 4951 5211 4994 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09884 4952 5818 4951 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09883 4950 5819 4952 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09882 7451 5815 4950 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09881 5241 4994 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09880 1316 1419 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09879 1468 1336 1316 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09878 7451 1337 1468 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09877 7451 1310 1308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09876 1307 1308 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09875 7451 1308 1307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09874 7451 1308 1307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09873 1307 1308 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09872 7451 1310 1311 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09871 1309 1311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09870 7451 1311 1309 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09869 7451 1311 1309 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09868 1309 1311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09867 7451 3246 2170 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09866 2169 2170 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09865 7451 2170 2169 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09864 7451 2170 2169 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09863 2169 2170 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09862 7451 3246 2247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09861 2246 2247 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09860 7451 2247 2246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09859 7451 2247 2246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09858 2246 2247 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09857 7451 3246 2248 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09856 2672 2248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09855 7451 2248 2672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09854 7451 2248 2672 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09853 2672 2248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09852 7451 3246 2178 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09851 2177 2178 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09850 7451 2178 2177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09849 7451 2178 2177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09848 2177 2178 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09847 7451 3246 2253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09846 2252 2253 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09845 7451 2253 2252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09844 7451 2253 2252 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09843 2252 2253 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09842 7451 3246 2254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09841 2533 2254 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09840 7451 2254 2533 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09839 7451 2254 2533 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09838 2533 2254 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09837 6970 7379 6950 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09836 6950 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09835 7451 7481 6970 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09834 6969 6970 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09833 7451 2111 918 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09832 7451 2602 919 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09831 918 919 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09830 2723 3911 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09829 7451 2860 2723 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09828 6109 6406 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09827 7451 7420 6108 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09826 7451 6323 6110 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09825 6126 6323 6109 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09824 6108 6110 6126 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09823 6107 6126 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09822 944 1550 926 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09821 926 1430 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09820 7451 1688 926 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09819 1336 944 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09818 925 1552 944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09817 926 1867 925 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09816 7451 3246 3164 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09815 3163 3164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09814 7451 3164 3163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09813 7451 3164 3163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09812 3163 3164 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09811 7451 3246 3236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09810 3235 3236 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09809 7451 3236 3235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09808 7451 3236 3235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09807 3235 3236 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09806 7451 3246 3237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09805 3581 3237 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09804 7451 3237 3581 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09803 7451 3237 3581 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09802 3581 3237 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09801 7451 3246 3169 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09800 3168 3169 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09799 7451 3169 3168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09798 7451 3169 3168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09797 3168 3169 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09796 7451 3246 3245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09795 3244 3245 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09794 7451 3245 3244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09793 7451 3245 3244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09792 3244 3245 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09791 7451 3246 3247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09790 3595 3247 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09789 7451 3247 3595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09788 7451 3247 3595 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09787 3595 3247 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09786 7451 3264 2188 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09785 2187 2188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09784 7451 2188 2187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09783 7451 2188 2187 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09782 2187 2188 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09781 7451 3304 3307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09780 3307 3411 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09779 7451 3412 3307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09778 3303 3307 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09777 4929 6534 4392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09776 4392 4815 4929 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09775 7451 4431 4392 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09774 7451 437 288 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09773 602 288 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09772 7451 288 602 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09771 7451 288 602 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09770 602 288 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09769 7451 602 395 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09768 5001 395 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09767 7451 395 5001 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09766 7451 395 5001 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09765 5001 395 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09764 7451 602 603 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09763 6133 603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09762 7451 603 6133 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09761 7451 603 6133 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09760 6133 603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09759 7451 3264 2259 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09758 2260 2259 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09757 7451 2259 2260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09756 7451 2259 2260 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09755 2260 2259 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09754 7451 3264 2262 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09753 2261 2262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09752 7451 2262 2261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09751 7451 2262 2261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09750 2261 2262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09749 7451 3264 2193 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09748 2192 2193 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09747 7451 2193 2192 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09746 7451 2193 2192 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09745 2192 2193 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09744 7451 3264 2266 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09743 2265 2266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09742 7451 2266 2265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09741 7451 2266 2265 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09740 2265 2266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09739 7451 3264 2267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09738 2553 2267 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09737 7451 2267 2553 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09736 7451 2267 2553 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09735 2553 2267 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09734 7451 3264 3177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09733 3176 3177 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09732 7451 3177 3176 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09731 7451 3177 3176 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09730 3176 3177 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09729 7451 3264 3254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09728 3253 3254 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09727 7451 3254 3253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09726 7451 3254 3253 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09725 3253 3254 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09724 7451 3264 3255 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09723 3466 3255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09722 7451 3255 3466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09721 7451 3255 3466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09720 3466 3255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09719 763 2222 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09718 7451 1851 763 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09717 762 763 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09716 1966 1965 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09715 7451 2157 1966 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09714 2091 1966 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09713 3450 3922 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09712 3513 3925 3450 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09711 7451 5138 3513 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09710 7451 6336 5903 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09709 5903 5905 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09708 5903 6477 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09707 7451 5902 5903 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09706 5904 5903 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09705 3926 5691 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09704 7451 5001 3926 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09703 3925 3926 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09702 7451 6979 6759 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09701 6759 6980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09700 7451 7464 6759 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09699 6757 6759 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09698 4096 4139 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09697 4094 4140 4134 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09696 7451 4933 4094 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09695 4140 4141 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09694 7451 4277 4141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09693 7451 4572 4139 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09692 4136 4140 4096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09691 4095 4141 4136 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09690 7451 4135 4095 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09689 4135 4136 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09688 4134 4141 4135 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09687 7451 4134 4933 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09686 4933 4134 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09685 6732 6965 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09684 4361 4933 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09683 2566 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09682 2589 2929 2566 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09681 7451 6035 2589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09680 7451 5691 3843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09679 3843 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09678 7451 5690 3843 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09677 3840 3843 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09676 6862 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09675 6899 7228 6862 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09674 7451 7475 6899 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09673 3724 3890 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09672 7173 7387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09671 7369 7480 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09670 6713 7045 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09669 7451 6991 6713 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09668 4807 5092 4825 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09667 4806 5716 4807 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09666 7451 4824 4806 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09665 6594 6682 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09664 7451 6593 6594 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09663 1204 1369 1175 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09662 1175 2255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09661 7451 4161 1204 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09660 1570 1204 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09659 1979 1631 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09658 7451 1581 1979 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09657 3186 3356 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09656 7451 3184 3186 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09655 3183 3186 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09654 6452 7267 6425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09653 6425 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09652 7451 7034 6425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09651 6451 6452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09650 6424 7032 6452 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09649 6425 7137 6424 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09648 1753 1898 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09647 7451 1688 1753 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09646 5166 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09645 5166 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09644 7451 5523 5166 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09643 7451 5690 5166 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09642 6286 6342 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09641 6608 6340 6286 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09640 7451 6341 6608 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09639 5090 5378 5091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09638 5088 6910 5090 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09637 5089 6981 5088 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09636 7451 5377 5089 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09635 5087 5091 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09634 4386 5138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09633 7451 5882 4385 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09632 7451 4912 4420 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09631 4419 4912 4386 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09630 4385 4420 4419 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09629 4416 4419 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09628 4201 5137 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09627 7451 6025 4200 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09626 7451 4912 4203 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09625 4202 4912 4201 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09624 4200 4203 4202 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09623 4475 4202 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09622 7451 4847 4849 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09621 4849 5071 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09620 7451 4848 4849 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09619 4846 4849 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09618 3082 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09617 7451 3226 3082 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09616 309 2708 325 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09615 324 1851 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09614 7451 324 309 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09613 3214 2171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09612 3214 2185 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09611 7451 4568 3214 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09610 4945 5365 4982 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09609 4983 5291 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09608 7451 4983 4945 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09607 4643 6030 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09606 4764 6029 4643 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09605 7451 5069 4764 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09604 7451 5521 5522 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09603 5522 7018 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09602 7451 5816 5522 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09601 5520 5522 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09600 2685 4000 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09599 2685 2684 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09598 7451 2687 2685 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09597 2649 2655 2651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09596 2650 2647 2649 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09595 7451 2648 2650 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09594 6165 2651 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09593 7451 6336 5993 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09592 5993 6112 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09591 7451 6576 5993 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09590 5992 5993 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09589 1417 1679 1418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09588 1418 1813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09587 7451 1684 1418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09586 1473 1417 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09585 1416 1680 1417 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09584 1418 1681 1416 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09583 774 828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09582 7451 908 774 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09581 1032 774 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09580 2523 3239 2524 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09579 2522 2521 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09578 7451 2522 2523 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09577 6958 7496 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09576 6957 7289 6958 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09575 7451 6981 6957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09574 3125 3214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09573 3145 3212 3125 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09572 7451 3879 3145 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09571 4147 4724 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09570 7451 5889 4147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09569 4224 4147 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09568 1993 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09567 2995 2541 1993 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09566 7451 2035 2995 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09565 7451 762 500 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09564 685 939 501 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09563 501 762 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09562 501 500 685 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09561 7451 499 501 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09560 499 939 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09559 7451 1051 734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09558 734 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09557 7451 2880 734 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09556 731 734 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09555 4163 4161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09554 7451 4376 4163 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09553 5172 4163 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09552 1313 2033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09551 7451 4600 1313 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09550 1312 1313 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09549 3887 3886 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09548 3880 3889 3881 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09547 7451 3879 3880 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09546 3889 3888 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09545 7451 4488 3888 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09544 7451 3884 3886 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09543 3885 3889 3887 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09542 3882 3888 3885 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09541 7451 3883 3882 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09540 3883 3885 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09539 3881 3888 3883 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09538 7451 3881 3879 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09537 3879 3881 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09536 7451 7164 4944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09535 4944 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09534 5364 4979 4944 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09533 4943 5275 5364 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09532 4944 5273 4943 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09531 3 16 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09530 1 17 11 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09529 7451 5125 1 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09528 17 18 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09527 7451 360 18 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09526 7451 5124 16 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09525 13 17 3 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09524 2 18 13 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09523 7451 12 2 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09522 12 13 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09521 11 18 12 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09520 7451 11 5125 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09519 5125 11 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09518 4384 4916 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09517 4415 4413 4384 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09516 4383 4411 4415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09515 7451 4412 4383 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09514 4410 4415 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09513 7451 4447 4235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09512 4235 4448 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09511 4235 4442 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09510 7451 4934 4235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09509 5842 4235 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09508 7004 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09507 7039 7228 7004 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09506 7451 7480 7039 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09505 6587 6852 6912 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09504 6653 7384 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09503 7451 6653 6587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09502 7451 4995 4931 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09501 4931 4996 4932 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09500 5273 4932 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09499 2986 4359 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09498 7451 3097 2986 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09497 5073 5072 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09496 7451 6944 5073 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09495 5071 5073 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09494 514 225 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09493 514 283 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09492 7451 518 514 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09491 641 1145 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09490 641 1029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09489 7451 640 641 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09488 7451 1809 641 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09487 7247 7309 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09486 7264 7416 7247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09485 7451 7420 7264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09484 6575 6576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09483 7451 7354 6575 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09482 6535 6575 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09481 7451 6534 4864 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09480 4864 5226 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09479 4864 4829 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09478 7451 4815 4864 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09477 5072 4864 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09476 2367 2418 2369 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09475 2369 2789 2368 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09474 2368 2505 2369 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09473 2367 2504 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09472 7451 2416 2367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09471 2369 2502 2367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09470 2366 2368 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09469 379 1082 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09468 7451 1688 379 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09467 378 379 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09466 7451 1976 1977 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09465 1977 2591 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09464 1977 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09463 7451 4376 1977 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09462 2542 1977 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09461 7451 4603 1839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09460 1839 4600 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09459 7451 7042 1839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09458 1838 1839 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09457 4528 4547 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09456 4526 4549 4541 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09455 7451 4975 4526 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09454 4549 4548 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09453 7451 4638 4548 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09452 7451 4641 4547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09451 4545 4549 4528 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09450 4527 4548 4545 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09449 7451 4543 4527 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09448 4543 4545 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09447 4541 4548 4543 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09446 7451 4541 4975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09445 4975 4541 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09444 7451 4448 4289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09443 4289 4441 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09442 4289 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09441 7451 4446 4289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09440 5718 4289 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09439 7451 1384 1298 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09438 1298 2392 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09437 1298 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09436 7451 2881 1298 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09435 1574 1298 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09434 4143 4069 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09433 7196 7453 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09432 7455 7454 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09431 4949 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09430 5082 5273 4949 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09429 7451 6035 5082 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09428 4243 4579 4274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09427 4244 5069 4243 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09426 7451 4774 4244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09425 4715 4274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09424 5367 5735 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09423 5366 5734 5367 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09422 7451 5815 5366 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09421 6323 7494 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09420 6770 7108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09419 2752 2889 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09418 7451 2751 2752 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09417 233 446 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09416 7451 3248 233 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09415 132 239 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09414 7451 4296 132 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09413 6308 6306 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09412 7451 6386 6308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09411 6310 6308 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09410 6825 6632 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09409 7451 6242 6825 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09408 4910 5369 4909 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09407 4909 4908 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09406 7451 5226 4910 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09405 5660 4910 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09404 6387 6389 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09403 7451 6386 6387 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09402 6633 6387 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09401 4681 4834 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09400 7451 6175 4680 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09399 7451 4912 4708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09398 4707 4912 4681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09397 4680 4708 4707 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09396 4705 4707 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09395 3757 5274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09394 7451 5887 3758 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09393 7451 4912 3788 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09392 3787 4912 3757 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09391 3758 3788 3787 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09390 4040 3787 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09389 275 1082 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09388 7451 1688 275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09387 3138 3403 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09386 7451 3137 3138 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09385 509 2696 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09384 7451 1851 509 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09383 2396 2540 2394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09382 2395 5841 2396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09381 2396 5840 2395 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09380 2394 2398 2396 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09379 2394 2536 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09378 7451 2684 2394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09377 7451 3074 2828 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09376 2829 3069 3633 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09375 2827 3070 2829 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09374 2828 3071 2827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09373 5540 5539 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09372 7451 5667 5540 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09371 5716 5904 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09370 7451 5891 5716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09369 7451 3351 3118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09368 3118 3119 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09367 7451 3266 3118 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09366 3181 3118 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09365 4683 5043 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09364 7451 6035 4682 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09363 7451 4912 4714 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09362 4712 4912 4683 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09361 4682 4714 4712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09360 4710 4712 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09359 2408 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09358 2662 2946 2408 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09357 7451 5216 2662 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09356 5844 7162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09355 5844 6332 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09354 7451 7042 5844 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09353 7451 1037 651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09352 651 2300 650 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09351 775 650 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09350 2087 2229 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09349 2659 2154 2087 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09348 7451 2164 2659 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09347 7451 4585 4587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09346 4587 4582 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09345 7451 4583 4587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09344 4581 4587 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09343 7451 6846 6723 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09342 6723 6770 6769 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09341 6768 6769 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09340 7451 558 365 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09339 6168 363 364 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09338 364 558 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09337 364 365 6168 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09336 7451 362 364 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09335 362 363 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09334 6131 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09333 6131 5718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09332 7451 4933 6131 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09331 7451 4934 6131 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09330 7451 1809 1269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09329 1269 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09328 2027 1339 1269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09327 1268 1266 2027 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09326 1269 1267 1268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09325 7451 1420 1421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09324 1421 1813 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09323 7451 1556 1421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09322 1419 1421 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09321 6712 6846 6711 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09320 6711 6770 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09319 7451 7354 6712 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09318 6710 6712 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09317 4487 4489 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09316 4482 4490 4484 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09315 7451 6035 4482 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09314 4490 4491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09313 7451 4488 4491 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09312 7451 4710 4489 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09311 4486 4490 4487 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09310 4485 4491 4486 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09309 7451 4483 4485 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09308 4483 4486 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09307 4484 4491 4483 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09306 7451 4484 6035 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09305 6035 4484 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09304 3423 3422 3966 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09303 7451 3820 3422 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09302 3424 3819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09301 3966 3820 3424 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09300 7451 3993 3423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09299 5687 5685 6394 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09298 5686 6333 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09297 7451 5686 5687 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09296 4343 4344 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09295 4338 4345 4339 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09294 7451 6175 4338 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09293 4345 4346 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09292 7451 4638 4346 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09291 7451 4705 4344 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09290 4342 4345 4343 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09289 4340 4346 4342 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09288 7451 4341 4340 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09287 4341 4342 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09286 4339 4346 4341 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09285 7451 4339 6175 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09284 6175 4339 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09283 7451 2171 1887 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09282 1887 2318 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09281 1887 2102 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09280 7451 4773 1887 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09279 4413 1887 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09278 7451 4377 1708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09277 1708 1707 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09276 1708 5173 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09275 7451 4376 1708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09274 1833 1708 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09273 305 1023 936 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09272 304 1022 305 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09271 7451 1021 304 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09270 7451 6553 6236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09269 6234 6629 6235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09268 6235 6553 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09267 6235 6236 6234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09266 7451 6233 6235 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09265 6233 6629 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09264 3741 3738 3740 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09263 3740 3739 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09262 7451 3736 3741 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09261 3737 3741 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09260 4701 6539 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09259 4701 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09258 7451 5826 4701 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09257 7451 7471 7362 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09256 7366 7475 7345 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09255 7345 7471 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09254 7345 7362 7366 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09253 7451 7363 7345 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09252 7363 7475 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09251 1997 2109 2183 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09250 1996 2042 1997 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09249 7451 2328 1996 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09248 3109 2954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09247 3109 2869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09246 7451 3179 3109 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09245 7451 2995 3109 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09244 6391 7494 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09243 6391 6967 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09242 7451 6968 6391 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09241 7451 325 82 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09240 225 186 83 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09239 83 325 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09238 83 82 225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09237 7451 81 83 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09236 81 186 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09235 7451 2602 920 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09234 921 1449 4442 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09233 922 1168 921 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09232 920 2111 922 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09231 3418 4985 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09230 3418 4368 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09229 7451 4367 3418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09228 7451 6408 3418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09227 1142 1332 1143 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09226 1143 1430 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09225 7451 3546 1143 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09224 1464 1142 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09223 1141 1333 1142 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09222 1143 1334 1141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09221 6554 7379 6524 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09220 6524 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09219 7451 6676 6554 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09218 6523 6554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09217 5569 5606 5607 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09216 5567 5818 5569 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09215 5568 5819 5567 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09214 7451 5815 5568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_09213 5828 5607 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09212 4299 5251 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09211 7451 4296 4299 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09210 4297 4299 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09209 1258 1144 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09208 7451 1342 1258 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09207 5696 5735 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09206 6681 5734 5696 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09205 7451 6315 6681 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09204 4925 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09203 4926 5273 4925 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09202 7451 6175 4926 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09201 3767 3819 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09200 7451 3993 3766 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09199 7451 3820 3823 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09198 3822 3820 3767 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09197 3766 3823 3822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09196 3817 3822 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09195 4724 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09194 4724 4603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09193 7451 4600 4724 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09192 7451 6333 4724 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09191 7451 7074 6729 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09190 6729 7452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09189 7451 7453 6729 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09188 6726 6729 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09187 1154 1866 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09186 1153 1270 1154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09185 1152 1342 1153 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09184 7451 1341 1152 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.22U AS=0.8372P AD=0.8372P PS=6.97U PD=6.97U 
Mtr_09183 5572 6770 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09182 5621 5620 5572 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09181 5573 6846 5621 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09180 7451 5619 5573 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09179 5685 5621 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09178 2646 2841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09177 7451 2836 2646 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09176 2645 2646 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09175 1901 2454 1844 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09174 1844 2816 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09173 7451 1899 1901 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09172 1898 1901 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09171 2656 3213 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09170 7451 2657 2656 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09169 2705 2656 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09168 7451 3033 3027 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09167 3027 3029 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09166 7451 3030 3027 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09165 3663 3027 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09164 4234 5172 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09163 7451 5171 4234 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09162 4603 4234 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09161 7451 1954 1676 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09160 3412 1858 1678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09159 1678 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09158 1678 1676 3412 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09157 7451 1677 1678 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09156 1677 1858 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09155 3898 3897 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09154 3891 3899 3893 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09153 7451 3890 3891 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09152 3899 3900 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09151 7451 4561 3900 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09150 7451 3895 3897 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09149 3896 3899 3898 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09148 3892 3900 3896 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09147 7451 3894 3892 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09146 3894 3896 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09145 3893 3900 3894 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09144 7451 3893 3890 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09143 3890 3893 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09142 6845 5001 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09141 3427 4148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09140 4805 4996 4823 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09139 4804 4822 4805 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09138 7451 7227 4804 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09137 3589 3593 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09136 3587 3594 3586 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09135 7451 3997 3587 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09134 3594 3596 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09133 7451 3595 3596 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_09132 7451 3592 3593 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09131 3590 3594 3589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09130 3591 3596 3590 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09129 7451 3588 3591 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09128 3588 3590 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09127 3586 3596 3588 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_09126 7451 3586 3997 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09125 3997 3586 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09124 3665 4156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09123 1709 1906 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09122 4593 5841 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09121 1572 1620 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09120 7451 1619 1572 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09119 980 978 933 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09118 933 1575 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09117 7451 1106 980 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09116 979 980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09115 4071 4360 4072 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09114 4072 4282 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09113 7451 6703 4071 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09112 4070 4071 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09111 7003 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09110 7103 7383 7003 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09109 7451 7452 7103 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09108 6750 6598 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09107 7451 6596 6750 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09106 3134 3135 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09105 7451 3644 3134 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09104 1549 1732 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09103 1641 1547 1549 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09102 7451 1548 1641 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09101 7283 4673 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09100 7451 4674 7283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09099 4757 4754 4758 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09098 4756 4755 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09097 7451 4756 4757 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09096 5081 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09095 5156 5273 5081 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09094 7451 6392 5156 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09093 6280 6323 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09092 6322 6406 6280 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09091 7451 7420 6322 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09090 887 5138 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09089 7451 3820 886 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09088 7451 6344 888 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09087 914 6344 887 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09086 886 888 914 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09085 915 914 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09084 657 5137 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09083 7451 4158 659 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09082 7451 6344 660 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09081 658 6344 657 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09080 659 660 658 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09079 656 658 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09078 811 5216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09077 7451 1168 810 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09076 7451 6344 870 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09075 869 6344 811 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09074 810 870 869 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09073 841 869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09072 1341 1700 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09071 1341 2718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09070 7451 1968 1341 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09069 7451 1688 1341 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09068 3735 3967 3731 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09067 5616 3732 3735 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09066 3735 3733 5616 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09065 3731 3734 3735 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09064 3731 3920 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09063 7451 4077 3731 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09062 4602 4603 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09061 7451 4600 4602 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09060 1148 1182 1147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09059 1147 1146 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09058 7451 1145 1148 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09057 1954 1148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09056 4821 4589 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09055 4821 4667 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09054 7451 4588 4821 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09053 2570 5055 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09052 7451 2602 2569 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09051 7451 6344 2607 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09050 2606 6344 2570 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09049 2569 2607 2606 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_09048 2603 2606 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09047 421 4161 1775 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09046 483 4376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09045 7451 483 421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09044 1299 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09043 1372 2541 1299 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09042 7451 1628 1372 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09041 1892 1896 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09040 1892 2104 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09039 7451 1893 1892 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09038 7451 6407 1892 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09037 5405 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09036 5451 6566 5405 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09035 7451 7454 5451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09034 1441 3820 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09033 1441 1976 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09032 7451 2392 1441 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09031 7451 4376 1441 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09030 5562 5885 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09029 5811 5884 5562 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09028 7451 6125 5811 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09027 1626 1624 1593 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09026 1593 1709 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09025 7451 4597 1626 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09024 1899 1626 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_09023 5857 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09022 6247 6394 5857 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09021 7451 5887 6247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09020 1229 1577 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09019 7451 3352 1229 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09018 2504 1229 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09017 7451 4368 4273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09016 4273 4367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09015 7451 4985 4273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09014 4566 4273 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09013 7451 6131 6130 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09012 6130 6708 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09011 7451 6533 6130 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09010 6705 6130 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09009 7451 4568 3716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09008 3716 4588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09007 7451 4569 3716 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_09006 4411 3716 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09005 7451 4069 3916 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09004 3916 4228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09003 7432 4378 3916 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09002 3915 4149 7432 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09001 3916 5909 3915 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_09000 5264 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08999 5460 5467 5264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08998 7451 7235 5460 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08997 3093 3094 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08996 3087 3095 3088 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08995 7451 3086 3087 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08994 3095 3096 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08993 7451 3571 3096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08992 7451 3092 3094 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08991 3091 3095 3093 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08990 3090 3096 3091 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08989 7451 3089 3090 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08988 3089 3091 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08987 3088 3096 3089 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08986 7451 3088 3086 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08985 3086 3088 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08984 6861 6894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08983 6976 6893 6861 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08982 7451 6892 6976 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08981 4196 6168 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08980 4195 6169 4196 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08979 7451 5069 4195 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08978 274 2134 273 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08977 273 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08976 7451 272 274 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08975 699 274 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08974 7451 7493 7332 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08973 7317 7494 7318 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08972 7318 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08971 7318 7332 7317 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08970 7451 7333 7318 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08969 7333 7494 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08968 6490 6611 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08967 7451 6490 6489 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08966 6488 6613 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08965 7451 6488 6421 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08964 6421 6489 6486 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08963 6486 6490 6420 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08962 6419 6491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08961 7451 6482 6491 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08960 6491 6482 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08959 6420 6483 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08958 6483 6486 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08957 7451 7500 6483 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08956 6482 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08955 6482 6489 6419 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08954 6483 6490 6482 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08953 3269 3293 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08952 3267 3294 3287 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08951 7451 3475 3267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08950 3294 3295 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08949 7451 3400 3295 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08948 7451 3476 3293 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08947 3290 3294 3269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08946 3268 3295 3290 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08945 7451 3289 3268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08944 3289 3290 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08943 3287 3295 3289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08942 7451 3287 3475 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08941 3475 3287 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08940 1980 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08939 2620 2541 1980 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08938 7451 1979 2620 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08937 4833 5045 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08936 4833 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08935 7451 5826 4833 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08934 6966 7016 6946 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08933 6946 7033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08932 7451 7034 6946 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08931 6944 6966 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08930 6945 7032 6966 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08929 6946 7307 6945 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08928 7451 3546 805 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08927 805 1430 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08926 827 900 805 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08925 804 823 827 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08924 805 824 804 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08923 467 3546 415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08922 7451 647 415 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08921 415 2016 467 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08920 464 467 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08919 1070 3545 1056 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08918 1056 2139 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08917 7451 1688 1070 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08916 1068 1070 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08915 7451 3927 3604 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08914 3605 4084 3660 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08913 3603 4006 3605 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08912 3604 3840 3603 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08911 5535 5677 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08910 7451 5534 5535 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08909 2435 2862 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08908 7451 2589 2435 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08907 1453 1883 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08906 7451 1699 1452 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08905 7451 3159 1487 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08904 1486 3159 1453 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08903 1452 1487 1486 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08902 1746 1486 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08901 2971 3266 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08900 2971 2825 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08899 7451 3119 2971 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08898 7451 3814 2971 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08897 7451 7164 4794 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08896 4794 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08895 4837 4834 4794 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08894 4793 5275 4837 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08893 4794 5273 4793 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08892 6008 7227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08891 6044 7228 6008 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08890 7451 7494 6044 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08889 3547 3549 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08888 3548 3545 3547 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08887 7451 3546 3548 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08886 7423 7477 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08885 7451 7480 7423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08884 7471 7423 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08883 6708 5000 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08882 6708 5718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08881 7451 5001 6708 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08880 306 893 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08879 363 455 306 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08878 7451 641 363 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08877 707 709 675 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08876 675 706 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08875 7451 1342 707 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08874 6030 707 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08873 7451 4728 4436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08872 4436 6133 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08871 7451 6333 4436 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08870 4996 4436 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08869 7451 6378 5732 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08868 5732 5728 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08867 7451 5729 5732 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08866 5727 5732 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08865 7451 7164 5058 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08864 5058 7286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08863 5056 5055 5058 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08862 5057 5275 5056 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08861 5058 5273 5057 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08860 5165 5166 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08859 7451 5451 5165 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08858 5306 5165 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08857 2466 2465 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08856 7451 2685 2466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08855 2463 2466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08854 7451 7489 7425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08853 7425 7481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08852 7425 7493 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08851 7451 7494 7425 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08850 7477 7425 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08849 107 108 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08848 103 109 102 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08847 7451 1906 103 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08846 109 110 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08845 7451 403 110 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08844 7451 132 108 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08843 105 109 107 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08842 106 110 105 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08841 7451 104 106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08840 104 105 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08839 102 110 104 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08838 7451 102 1906 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08837 1906 102 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08836 4768 5376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08835 4921 5273 4768 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08834 7451 6025 4921 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08833 1084 1430 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08832 7451 1466 1084 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08831 3545 1084 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08830 3485 3484 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08829 7451 3483 3485 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08828 3482 3485 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08827 1770 2395 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08826 7451 1767 1770 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08825 1768 1770 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08824 1323 2255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08823 1568 1363 1323 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08822 7451 1449 1568 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08821 795 1112 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08820 7451 1111 795 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08819 1047 795 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08818 7451 7105 7106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08817 7106 7103 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08816 7451 7156 7106 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08815 7104 7106 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08814 7451 6979 6127 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08813 6127 6980 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08812 7451 7466 6127 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08811 6111 6127 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08810 420 918 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08809 729 481 420 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08808 7451 3427 729 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08807 7451 3727 3728 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08806 3728 4228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08805 5835 3819 3728 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08804 3726 4149 5835 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08803 3728 5909 3726 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08802 7451 4081 244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08801 244 4437 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08800 7451 5001 244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08799 242 244 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08798 7451 1736 208 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08797 1633 890 197 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08796 197 1736 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08795 197 208 1633 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08794 7451 206 197 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08793 206 890 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08792 5112 5147 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08791 5110 5148 5141 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08790 7451 5833 5110 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08789 5148 5149 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08788 7451 5518 5149 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08787 7451 5229 5147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08786 5144 5148 5112 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08785 5111 5149 5144 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08784 7451 5143 5111 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08783 5143 5144 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08782 5141 5149 5143 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08781 7451 5141 5833 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08780 5833 5141 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08779 2255 2602 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08778 2103 4161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08777 5000 4934 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08776 171 1022 172 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08775 172 1021 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08774 7451 1023 171 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08773 937 171 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08772 7451 1435 1424 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08771 1424 1768 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08770 1422 1556 1424 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08769 1423 1682 1422 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08768 1424 1479 1423 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08767 4296 1508 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08766 7451 7162 4296 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08765 7451 6869 6623 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08764 6625 6732 6577 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08763 6577 6869 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08762 6577 6623 6625 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08761 7451 6624 6577 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08760 6624 6732 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08759 6466 6697 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08758 7451 6464 6466 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08757 5329 7390 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08756 6135 6652 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08755 4822 4780 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08754 7451 4781 4822 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08753 6690 6032 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08752 7451 6033 6690 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08751 5654 5653 5668 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08750 5652 5818 5654 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08749 5651 5819 5652 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08748 7451 5815 5651 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.25U AS=0.585P AD=0.585P PS=5.02U PD=5.02U 
Mtr_08747 5669 5668 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08746 829 828 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08745 7451 908 829 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08744 7110 7109 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08743 7451 7108 7110 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08742 3143 3079 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08741 3143 3080 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08740 7451 3482 3143 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08739 1567 1883 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08738 7451 1699 1567 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08737 4820 4773 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08736 4820 4568 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08735 7451 4569 4820 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08734 4726 7162 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08733 4726 2033 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08732 7451 4600 4726 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08731 2418 2228 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08730 2418 4694 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08729 7451 2524 2418 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08728 6004 6030 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08727 6033 6029 6004 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08726 7451 6315 6033 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08725 5069 4367 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08724 5069 5085 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08723 7451 4368 5069 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08722 7451 4985 5069 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08721 1998 2543 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08720 2256 2541 1998 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08719 7451 2179 2256 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08718 7451 2988 2957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08717 2957 2958 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08716 7451 2956 2957 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08715 6046 2957 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08714 5300 5274 5121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08713 5121 5832 5300 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08712 7451 5153 5121 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08711 2375 3418 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08710 2657 2929 2375 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08709 7451 6392 2657 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08708 4083 4161 4447 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08707 4082 4158 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08706 7451 4082 4083 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08705 6058 6773 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08704 6058 6535 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08703 7451 6114 6058 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08702 7451 6056 6058 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08701 4657 4659 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08700 4653 4661 4654 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08699 7451 5454 4653 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08698 4661 4662 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08697 7451 4660 4662 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08696 7451 4779 4659 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08695 4658 4661 4657 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08694 4656 4662 4658 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08693 7451 4655 4656 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08692 4655 4658 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08691 4654 4662 4655 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08690 7451 4654 5454 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08689 5454 4654 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08688 2136 3131 2122 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08687 2122 2286 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08686 7451 2133 2136 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08685 2134 2136 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08684 923 936 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08683 3469 937 923 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08682 7451 1342 3469 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08681 2981 3501 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08680 3719 4669 2981 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08679 7451 3226 3719 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08678 3645 4431 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08677 3226 4991 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08676 889 2095 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08675 890 3545 889 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08674 7451 1688 890 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08673 1065 3545 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08672 3917 2027 1065 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08671 7451 2029 3917 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08670 3646 4718 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08669 3012 4424 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08668 4378 4937 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08667 7451 1236 794 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08666 794 1441 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08665 7451 844 794 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08664 978 794 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08663 537 1052 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08662 7451 1775 537 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08661 536 537 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08660 5508 6894 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08659 5581 5902 5508 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08658 7451 5507 5581 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08657 546 588 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08656 544 587 580 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08655 7451 579 544 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08654 587 589 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08653 7451 788 589 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08652 7451 584 588 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08651 585 587 546 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08650 545 589 585 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08649 7451 582 545 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08648 582 585 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08647 580 589 582 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08646 7451 580 579 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08645 579 580 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08644 3404 4695 3405 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08643 3405 3481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08642 7451 3484 3404 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08641 3403 3404 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08640 1071 1337 1062 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08639 1062 1952 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08638 7451 1548 1062 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08637 1074 1071 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08636 1061 1419 1071 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08635 1062 1336 1061 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08634 4041 4043 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08633 4036 4045 4037 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08632 7451 5887 4036 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08631 4045 4044 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08630 7451 4638 4044 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08629 7451 4040 4043 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08628 4042 4045 4041 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08627 4038 4044 4042 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08626 7451 4039 4038 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08625 4039 4042 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08624 4037 4044 4039 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08623 7451 4037 5887 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08622 5887 4037 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08621 298 403 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08620 7451 298 297 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08619 296 295 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08618 7451 296 293 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08617 293 297 294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08616 294 298 291 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08615 289 4376 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08614 7451 290 4376 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08613 4376 290 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08612 291 292 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08611 292 294 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08610 7451 7500 292 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08609 290 7500 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08608 290 297 289 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08607 292 298 290 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.02U AS=0.5252P AD=0.5252P PS=4.57U PD=4.57U 
Mtr_08606 6142 6393 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08605 6318 6394 6142 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08604 7451 6175 6318 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08603 7451 195 196 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08602 196 242 405 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08601 4664 4821 4777 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08600 4663 4819 4664 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08599 7451 4820 4663 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08598 2799 2854 2803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08597 2803 2800 2802 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08596 2802 2801 2803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08595 2799 2991 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08594 7451 2995 2799 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08593 2803 4410 2799 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08592 2798 2802 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08591 3918 3917 3919 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08590 3919 5889 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08589 7451 4825 3918 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08588 4075 3918 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08587 5498 5350 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08586 5498 5351 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08585 7451 5826 5498 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08584 942 2222 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08583 7451 1851 942 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08582 1554 1867 1553 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08581 1553 1552 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08580 7451 1550 1554 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08579 1551 1554 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08578 7451 7264 6879 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08577 6879 6878 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08576 7451 6947 6879 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08575 6876 6879 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08574 5302 5300 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08573 7451 5299 5302 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08572 5438 5302 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08571 2793 3481 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08570 2792 4695 2793 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08569 7451 3077 2792 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08568 6762 7104 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08567 7451 6761 6762 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08566 7451 5312 4223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08565 4222 4223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08564 7451 4223 4222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08563 7451 4223 4222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08562 4222 4223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08561 7451 5312 4276 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08560 4275 4276 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08559 7451 4276 4275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08558 7451 4276 4275 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08557 4275 4276 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08556 7451 5312 4278 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08555 4277 4278 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08554 7451 4278 4277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08553 7451 4278 4277 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08552 4277 4278 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08551 7451 5312 4227 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08550 4226 4227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08549 7451 4227 4226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08548 7451 4227 4226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08547 4226 4227 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08546 7451 5312 4284 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08545 4283 4284 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08544 7451 4284 4283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08543 7451 4284 4283 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08542 4283 4284 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08541 7451 5312 4285 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08540 4660 4285 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08539 7451 4285 4660 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08538 7451 4285 4660 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08537 4660 4285 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08536 7451 5312 5240 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08535 5239 5240 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08534 7451 5240 5239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08533 7451 5240 5239 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08532 5239 5240 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08531 314 1681 300 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08530 300 1680 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08529 7451 1679 314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08528 312 314 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08527 2008 1809 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08526 2008 1954 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08525 7451 1810 2008 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08524 2618 3431 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08523 2618 4524 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08522 7451 2620 2618 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08521 7451 2823 2618 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08520 270 1021 455 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08519 269 462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08518 7451 269 270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08517 2974 3137 2975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08516 2975 2991 2992 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08515 2992 2995 2975 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08514 2974 3082 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08513 7451 3701 2974 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08512 2975 3403 2974 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08511 3406 2992 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08510 1345 1341 1318 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08509 1318 1340 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08508 7451 1342 1318 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08507 1339 1345 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08506 1317 1551 1345 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08505 1318 1741 1317 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08504 7451 5312 5304 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08503 5303 5304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08502 7451 5304 5303 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08501 7451 5304 5303 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08500 5303 5304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08499 7451 5312 5305 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08498 5531 5305 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08497 7451 5305 5531 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08496 7451 5305 5531 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08495 5531 5305 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08494 7451 5312 5246 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08493 5245 5246 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08492 7451 5246 5245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08491 7451 5246 5245 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08490 5245 5246 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08489 7451 5312 5311 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08488 5310 5311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08487 7451 5311 5310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08486 7451 5311 5310 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08485 5310 5311 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08484 7451 5312 5313 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08483 5449 5313 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08482 7451 5313 5449 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08481 7451 5313 5449 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08480 5449 5313 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08479 7451 5327 4233 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08478 4232 4233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08477 7451 4233 4232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08476 7451 4233 4232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08475 4232 4233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08474 7451 5327 4293 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08473 4292 4293 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08472 7451 4293 4292 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08471 7451 4293 4292 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08470 4292 4293 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08469 7451 5327 4295 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08468 4294 4295 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08467 7451 4295 4294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08466 7451 4295 4294 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08465 4294 4295 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08464 1738 1876 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08463 7451 1851 1738 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08462 1736 1738 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08461 7451 3160 2952 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08460 2952 3303 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08459 2952 3159 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08458 7451 3326 2952 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08457 2951 2952 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08456 6138 6234 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08455 6162 6160 6138 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08454 7451 7420 6162 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08453 2839 3128 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08452 7451 2836 2839 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08451 2837 2839 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08450 6430 6565 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08449 6473 6566 6430 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08448 7451 7335 6473 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08447 7451 5327 4237 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08446 4236 4237 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08445 7451 4237 4236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08444 7451 4237 4236 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08443 4236 4237 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08442 7451 5327 4304 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08441 4303 4304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08440 7451 4304 4303 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08439 7451 4304 4303 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08438 4303 4304 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08437 7451 5327 4306 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08436 4305 4306 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08435 7451 4306 4305 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08434 7451 4306 4305 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08433 4305 4306 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08432 7451 5327 5248 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08431 5247 5248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08430 7451 5248 5247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08429 7451 5248 5247 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08428 5247 5248 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08427 7451 5327 5318 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08426 5317 5318 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08425 7451 5318 5317 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08424 7451 5318 5317 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08423 5317 5318 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08422 7451 5327 5320 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08421 5319 5320 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08420 7451 5320 5319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08419 7451 5320 5319 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08418 5319 5320 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08417 7451 5327 5255 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08416 5254 5255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08415 7451 5255 5254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08414 7451 5255 5254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08413 5254 5255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08412 2509 2856 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08411 7451 2657 2509 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08410 2846 2509 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08409 341 399 303 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08408 303 340 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08407 7451 5619 341 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08406 1109 341 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08405 1606 3546 1586 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08404 1586 1883 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08403 7451 1851 1586 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08402 1605 1606 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08401 1585 1823 1606 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08400 1586 3545 1585 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08399 7451 1876 1878 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08398 1878 2424 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08397 7451 2220 1878 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08396 2093 1878 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08395 7451 7413 7324 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08394 7307 7462 7308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08393 7308 7413 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08392 7308 7324 7307 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08391 7451 7325 7308 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08390 7325 7462 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08389 7451 775 575 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08388 575 1155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08387 7451 1688 575 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08386 653 575 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08385 7451 2718 1036 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08384 1036 1968 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08383 7451 1700 1036 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08382 1430 1036 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08381 2030 2029 1992 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08380 1992 5889 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08379 7451 4568 1992 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08378 2820 2030 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08377 1991 3545 2030 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08376 1992 2027 1991 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08375 7451 5327 5326 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08374 5325 5326 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08373 7451 5326 5325 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08372 7451 5326 5325 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08371 5325 5326 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08370 7451 5327 5328 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08369 5554 5328 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08368 7451 5328 5554 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08367 7451 5328 5554 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08366 5554 5328 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08365 7451 7224 6178 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08364 6177 6178 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08363 7451 6178 6177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08362 7451 6178 6177 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08361 6177 6178 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08360 7451 7224 6250 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08359 6249 6250 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08358 7451 6250 6249 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08357 7451 6250 6249 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08356 6249 6250 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08355 7451 7224 6251 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08354 6693 6251 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08353 7451 6251 6693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08352 7451 6251 6693 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08351 6693 6251 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08350 7451 7224 6184 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08349 6183 6184 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08348 7451 6184 6183 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08347 7451 6184 6183 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08346 6183 6184 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08345 7451 7224 6255 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08344 6254 6255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08343 7451 6255 6254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08342 7451 6255 6254 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08341 6254 6255 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08340 7451 7224 6257 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08339 6256 6257 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08338 7451 6257 6256 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08337 7451 6257 6256 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08336 6256 6257 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08335 3939 3987 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08334 3937 3986 3984 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08333 7451 4215 3937 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08332 3986 3988 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08331 7451 4277 3988 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08330 7451 4216 3987 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08329 3961 3986 3939 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08328 3938 3988 3961 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08327 7451 3960 3938 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08326 3960 3961 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08325 3984 3988 3960 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08324 7451 3984 4215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08323 4215 3984 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08322 517 3081 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08321 518 1085 517 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08320 7451 775 518 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08319 6549 4702 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08318 7451 4249 6549 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08317 5215 5214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08316 7451 6672 5215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08315 5095 5249 5097 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08314 5096 5688 5095 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08313 7451 5378 5096 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08312 4512 5832 4514 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08311 4513 4827 4512 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08310 7451 4511 4513 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08309 7451 7224 7148 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08308 7147 7148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08307 7451 7148 7147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08306 7451 7148 7147 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08305 7147 7148 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08304 7451 7224 7214 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08303 7213 7214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08302 7451 7214 7213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08301 7451 7214 7213 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08300 7213 7214 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08299 7451 7224 7216 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08298 7215 7216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08297 7451 7216 7215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08296 7451 7216 7215 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08295 7215 7216 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08294 7451 7224 7155 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08293 7154 7155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08292 7451 7155 7154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08291 7451 7155 7154 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08290 7154 7155 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08289 7451 7224 7223 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08288 7222 7223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08287 7451 7223 7222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08286 7451 7223 7222 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08285 7222 7223 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08284 7451 7224 7226 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08283 7225 7226 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08282 7451 7226 7225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08281 7451 7226 7225 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08280 7225 7226 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08279 7451 7474 7327 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08278 7313 7466 7314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08277 7314 7474 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08276 7314 7327 7313 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08275 7451 7328 7314 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08274 7328 7466 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08273 655 653 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08272 910 654 655 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08271 7451 833 910 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08270 7354 7353 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08269 7451 7384 7354 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08268 3120 6340 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08267 7451 3516 3120 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08266 7451 7240 6192 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08265 6191 6192 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08264 7451 6192 6191 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08263 7451 6192 6191 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08262 6191 6192 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08261 908 907 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08260 7451 1341 908 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08259 4368 7042 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08258 4368 1292 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08257 7451 4600 4368 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08256 6722 7334 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08255 6764 7383 6722 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08254 7451 6965 6764 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08253 5803 7452 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08252 5803 6156 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08251 7451 6968 5803 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08250 7451 7240 6262 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08249 6261 6262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08248 7451 6262 6261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08247 7451 6262 6261 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08246 6261 6262 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08245 7451 7240 6264 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08244 6263 6264 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08243 7451 6264 6263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08242 7451 6264 6263 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08241 6263 6264 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08240 7451 7240 6200 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08239 6199 6200 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08238 7451 6200 6199 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08237 7451 6200 6199 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08236 6199 6200 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08235 7451 7240 6269 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08234 6268 6269 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08233 7451 6269 6268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08232 7451 6269 6268 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08231 6268 6269 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08230 7248 7491 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08229 7267 7379 7248 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08228 7451 7464 7267 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08227 2131 3837 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08226 2190 2467 2131 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08225 2130 2337 2190 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08224 7451 2338 2130 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08223 2189 2190 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08222 5889 6333 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08221 5889 5842 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08220 7451 5841 5889 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08219 2026 2946 1990 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08218 1990 2945 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08217 7451 5138 2026 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08216 2099 2026 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.32U AS=0.6032P AD=0.6032P PS=5.17U PD=5.17U 
Mtr_08215 7244 7513 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08214 7440 7243 7244 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08213 7451 7242 7440 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08212 7451 7240 6270 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08211 6611 6270 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08210 7451 6270 6611 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08209 7451 6270 6611 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08208 6611 6270 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08207 7451 7240 7161 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08206 7160 7161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08205 7451 7161 7160 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08204 7451 7161 7160 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08203 7160 7161 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08202 7451 7240 7231 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08201 7230 7231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08200 7451 7231 7230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08199 7451 7231 7230 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08198 7230 7231 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08197 7451 7240 7233 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08196 7232 7233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08195 7451 7233 7232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08194 7451 7233 7232 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08193 7232 7233 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08192 4598 6576 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08191 7451 4597 4598 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08190 5459 4598 7451 7451 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.92U AS=0.7592P AD=0.7592P PS=6.37U PD=6.37U 
Mtr_08189 7514 7240 7171 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08188 7170 7171 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08187 7514 7171 7170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08186 7514 7171 7170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08185 7170 7171 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08184 7514 1170 4446 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08183 1170 1168 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08182 4446 1449 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08181 2049 2412 2050 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08180 2050 2645 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08179 3067 2922 2049 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08178 7514 1021 357 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08177 7514 1022 357 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08176 357 1023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08175 1020 357 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08174 5671 6316 5603 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08173 5603 6314 5671 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08172 7514 5815 5603 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08171 7514 7240 7239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08170 7238 7239 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08169 7514 7239 7238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08168 7514 7239 7238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08167 7238 7239 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08166 7514 7240 7241 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08165 7508 7241 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08164 7514 7241 7508 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08163 7514 7241 7508 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08162 7508 7241 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08161 7514 6771 4776 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08160 5312 4776 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08159 7514 4776 5312 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08158 7514 4776 5312 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08157 5312 4776 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08156 6596 6316 6317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08155 6317 6314 6596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08154 7514 6315 6317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08153 3100 3105 3101 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08152 3051 3107 3100 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08151 4424 3100 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08150 7514 3100 4424 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08149 3054 3106 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08148 7514 3324 3106 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08147 3105 3107 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08146 7514 3581 3107 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08145 3052 3104 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08144 3101 5100 3052 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08143 3104 3107 3054 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08142 3053 3105 3104 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08141 7514 3101 3053 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08140 7514 4424 3050 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08139 3050 5100 3051 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08138 7514 6771 4788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08137 5327 4788 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08136 7514 4788 5327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08135 7514 4788 5327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08134 5327 4788 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08133 7514 6771 6756 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08132 7224 6756 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08131 7514 6756 7224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08130 7514 6756 7224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08129 7224 6756 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08128 7514 6771 6772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08127 7240 6772 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08126 7514 6772 7240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08125 7514 6772 7240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08124 7240 6772 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08123 7514 4588 1617 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08122 1617 1832 1654 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08121 1653 1654 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08120 7514 6907 6909 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08119 6909 7044 6908 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08118 6906 6908 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08117 2661 3149 2628 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08116 2628 4695 2661 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08115 7514 2856 2628 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08114 7514 7384 7386 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08113 7386 7391 7385 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08112 7383 7385 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08111 7514 5752 1739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08110 2712 1739 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08109 7514 1739 2712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08108 7514 1739 2712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08107 2712 1739 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08106 7514 5752 1762 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08105 2746 1762 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08104 7514 1762 2746 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08103 7514 1762 2746 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08102 2746 1762 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08101 716 1040 715 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08100 715 1041 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08099 714 4588 716 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08098 832 713 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_08097 713 4589 714 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08096 47 72 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_08095 45 74 66 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08094 7514 4104 45 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08093 7514 368 74 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_08092 73 74 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_08091 7514 4103 72 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_08090 68 69 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08089 7514 68 46 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08088 66 73 68 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08087 4104 66 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08086 7514 66 4104 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08085 46 73 69 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08084 69 74 47 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_08083 4889 5171 4890 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08082 4890 5172 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08081 4888 5173 4889 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08080 6566 4935 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_08079 4935 7042 4888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08078 725 1168 726 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08077 726 4161 727 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08076 7514 4376 725 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08075 1292 727 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_08074 5667 5734 5632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08073 5632 5735 5667 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08072 7514 6125 5632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08071 3524 3562 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08070 6314 3563 3524 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08069 3382 3487 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08068 3804 3409 3382 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08067 2293 3023 2295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08066 2294 2292 2293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08065 2295 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08064 2652 2293 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08063 7514 2583 2294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08062 2294 3549 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08061 7514 6386 6352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08060 6352 6384 6385 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08059 6878 6385 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08058 7514 4703 4702 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08057 4703 4701 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08056 4702 5215 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08055 4977 5826 4976 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08054 4976 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08053 4978 4975 4977 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08052 638 2576 614 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08051 613 3546 638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08050 614 1851 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08049 1679 638 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08048 7514 3549 613 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08047 613 3545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_08046 7514 5287 5420 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08045 5287 5286 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08044 5420 5417 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08043 4612 5826 4611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08042 4611 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08041 4847 4642 4612 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08040 2775 3170 2774 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08039 2774 3655 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08038 3343 5138 2775 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08037 7514 4411 4256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_08036 4256 4255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_08035 4254 4257 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08034 4256 4413 4257 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_08033 4257 4841 4256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_08032 2417 2416 2419 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08031 2419 2418 2420 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08030 2420 2789 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08029 2415 2504 2419 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08028 7514 2424 2415 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08027 7514 2502 2417 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08026 2648 2419 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08025 7326 7491 7292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08024 7292 7379 7326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08023 7514 7464 7292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08022 7309 7326 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08021 7514 2956 2317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08020 2317 2676 2316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08019 2315 2316 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08018 2228 3418 2015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08017 2015 2929 2228 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08016 7514 6175 2015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08015 7514 2288 1789 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08014 1789 2023 1818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08013 1821 1818 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08012 7514 2958 2903 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08011 2903 2988 2959 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08010 3030 2959 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_08009 5464 5459 5465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08008 5465 5460 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08007 5462 6405 5464 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08006 5905 5463 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_08005 5463 5461 5462 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08004 5893 5891 5894 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08003 5894 5992 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08002 5892 5902 5893 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_08001 6156 5890 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_08000 5890 5889 5892 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07999 2496 2552 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07998 2494 2554 2546 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07997 7514 7108 2494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07996 7514 2553 2554 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07995 2551 2554 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07994 7514 2752 2552 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07993 2547 2550 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07992 7514 2547 2495 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07991 2546 2551 2547 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07990 7108 2546 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07989 7514 2546 7108 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07988 2495 2551 2550 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07987 2550 2554 2496 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07986 7514 7108 4626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07985 4626 5691 4678 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07984 4679 4678 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07983 7236 7387 7185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07982 7185 7512 7236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07981 7514 7235 7185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07980 7037 7033 7036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07979 7035 7101 7037 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07978 7036 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07977 7031 7037 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07976 7514 7032 7035 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07975 7035 7317 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07974 6288 6292 6291 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07973 7514 7452 6288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07972 6290 6518 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07971 6291 6289 6290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07970 7514 6518 6292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07969 6289 7452 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07968 5534 6030 5298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07967 5298 6029 5534 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07966 7514 5815 5298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07965 1875 1871 1874 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07964 1874 1872 1873 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07963 7514 2798 1875 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07962 2018 1873 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07961 1498 1620 1499 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07960 1497 1834 1498 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07959 1499 1619 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07958 1496 1498 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07957 7514 3425 1497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07956 1497 1631 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07955 3866 5001 3867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07954 3867 5842 3928 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07953 7514 5690 3866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07952 3927 3928 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07951 877 1435 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07950 903 1768 877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07949 876 902 903 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07948 7514 899 876 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07947 876 900 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07946 4748 4837 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07945 4752 6009 4748 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07944 2736 2748 2737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07943 2737 2741 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07942 2735 5093 2736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07941 2733 2734 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07940 2734 4732 2735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07939 5085 6566 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07938 7514 6565 5085 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07937 4111 4758 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07936 4966 4195 4111 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07935 4704 5218 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07934 4754 6150 4704 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07933 777 960 623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07932 623 832 777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07931 7514 2592 623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07930 1123 1605 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07929 1340 1426 1123 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07928 3694 5623 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07927 6342 6333 3694 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07926 2910 3259 2911 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07925 2911 2972 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07924 2973 2971 2910 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07923 7514 6030 3713 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07922 3713 3957 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07921 7514 3958 3713 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07920 4826 5097 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07919 4827 4829 4826 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07918 149 179 563 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07917 7514 509 149 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07916 150 181 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07915 563 180 150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07914 7514 181 179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07913 180 509 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07912 2912 3135 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07911 2931 3500 2912 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07910 5266 5987 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07909 5267 5664 5266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07908 939 2139 940 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07907 940 3545 939 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07906 7514 1688 940 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07905 7514 6907 6478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07904 6478 6843 6479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07903 6477 6479 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07902 6157 6968 6159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07901 6159 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07900 6158 7453 6157 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07899 456 502 3409 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07898 7514 691 456 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07897 457 894 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07896 3409 503 457 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07895 7514 894 502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07894 503 691 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07893 1414 2095 1389 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07892 1389 3545 1414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07891 7514 1688 1389 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07890 1413 1414 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07889 5756 5844 5759 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07888 5759 5913 5758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07887 7514 6267 5756 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07886 5757 5758 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07885 2062 2171 2061 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07884 2061 2318 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07883 2060 2102 2062 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07882 2925 4773 2060 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07881 2883 4446 2882 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07880 2882 2880 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07879 4674 2881 2883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07878 4848 5275 4736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07877 4736 5273 4848 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07876 7514 5043 4736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07875 1820 1821 1790 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07874 1790 1823 1820 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07873 7514 2154 1790 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07872 1819 1820 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07871 3565 3572 3566 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07870 3527 3574 3565 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07869 4991 3565 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07868 7514 3565 4991 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07867 3529 3573 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07866 7514 3568 3573 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07865 3572 3574 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07864 7514 3571 3574 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07863 3526 3570 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07862 3566 7500 3526 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07861 3570 3574 3529 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07860 3528 3572 3570 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07859 7514 3566 3528 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07858 7514 4991 3525 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07857 3525 7500 3527 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07856 2413 3129 2414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07855 2414 4695 2413 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07854 7514 3128 2414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07853 2412 2413 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07852 5740 5743 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07851 5712 5744 5739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07850 7514 6187 5712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07849 7514 6693 5744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07848 5742 5744 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07847 7514 5741 5743 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07846 5713 5714 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07845 7514 5713 5715 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07844 5739 5742 5713 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07843 6187 5739 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07842 7514 5739 6187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07841 5715 5742 5714 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07840 5714 5744 5740 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07839 7514 3546 154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07838 154 2016 187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07837 186 187 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07836 688 1145 690 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07835 690 1029 689 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07834 7514 1809 688 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07833 1021 689 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07832 1435 2174 1404 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07831 1404 1837 1435 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07830 7514 6333 1404 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07829 7514 1384 1387 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07828 1387 1385 1386 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07827 2033 1386 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07826 7025 7022 7024 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07825 7514 7481 7025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07824 7026 7095 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07823 7024 7023 7026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07822 7514 7095 7022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07821 7023 7481 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07820 2208 2880 2209 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07819 2209 2263 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07818 2207 4446 2208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07817 2540 2264 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07816 2264 2881 2207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07815 7514 2044 2398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07814 2044 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07813 2398 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07812 6569 6565 6329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07811 6329 6566 6569 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07810 7514 6965 6329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07809 750 786 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07808 748 789 780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07807 7514 4161 748 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07806 7514 788 789 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07805 787 789 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07804 7514 785 786 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07803 781 784 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07802 7514 781 749 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07801 780 787 781 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07800 4161 780 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07799 7514 780 4161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07798 749 787 784 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07797 784 789 750 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07796 1726 1893 1725 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07795 1725 2104 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07794 1724 1896 1726 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07793 1825 1756 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07792 1756 6407 1724 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07791 137 135 266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07790 7514 3548 137 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07789 138 1852 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07788 266 136 138 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07787 7514 1852 135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07786 136 3548 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07785 7514 3997 3371 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07784 3371 4577 3419 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07783 7514 4577 3392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07782 3419 3392 3372 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07781 3592 3419 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07780 3372 3389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07779 6377 7491 6348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07778 6348 7379 6377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07777 7514 7335 6348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07776 6375 6377 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07775 7514 4933 4573 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07774 4573 4577 4576 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07773 7514 4577 4578 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07772 4576 4578 4575 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07771 4572 4576 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07770 4575 4574 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07769 7514 3890 3640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07768 3640 4577 3641 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07767 7514 4577 3642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07766 3641 3642 3643 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07765 3895 3641 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07764 3643 3870 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07763 7514 4215 4181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07762 4181 4577 4220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07761 7514 4577 4221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07760 4220 4221 4182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07759 4216 4220 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07758 4182 4217 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07757 2498 2537 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07756 2727 7162 2498 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07755 5772 5810 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07754 5812 5811 5772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07753 4003 6133 4002 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07752 4002 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07751 4001 4000 4003 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07750 5461 6333 4001 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07749 7514 4820 4865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07748 7514 4819 4865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07747 4865 4821 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07746 5815 4865 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07745 2526 2531 2527 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07744 2487 2534 2526 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07743 3819 2526 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07742 7514 2526 3819 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07741 2490 2532 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07740 7514 2866 2532 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07739 2531 2534 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07738 7514 2533 2534 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07737 2488 2529 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07736 2527 7500 2488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07735 2529 2534 2490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07734 2489 2531 2529 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07733 7514 2527 2489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07732 7514 3819 2486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07731 2486 7500 2487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07730 6982 6987 6984 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07729 6930 6983 6982 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07728 6991 6982 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07727 7514 6982 6991 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07726 6933 6986 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07725 7514 6988 6986 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07724 6987 6983 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07723 7514 7508 6983 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07722 6931 6985 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07721 6984 7500 6931 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07720 6985 6983 6933 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07719 6932 6987 6985 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07718 7514 6984 6932 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07717 7514 6991 6929 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07716 6929 7500 6930 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07715 7422 7419 7396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07714 7396 7470 7422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07713 7514 7420 7396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07712 4570 4568 4571 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07711 4571 5369 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07710 5275 4569 4570 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07709 3542 3817 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07708 3734 3837 3542 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07707 1870 3000 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07706 1867 1869 1870 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07705 1868 3546 1867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07704 7514 2095 1868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07703 1868 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07702 7514 963 838 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07701 838 875 863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07700 7514 875 864 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07699 863 864 837 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07698 968 863 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07697 837 3917 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07696 1155 2435 1125 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07695 1125 2853 1155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07694 7514 2133 1125 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07693 5323 6061 5322 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07692 5322 6652 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07691 5324 7390 5323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07690 5466 7388 5324 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07689 2301 3645 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07688 2300 3135 2301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07687 2299 2926 2300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07686 7514 6035 2299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07685 2298 2925 2300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07684 7514 5043 2298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07683 778 3081 488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07682 488 1085 778 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07681 7514 831 488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07680 7514 3409 3301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07679 3301 3487 3302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07678 3300 3302 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07677 7514 4411 3007 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07676 3007 3005 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07675 3004 3006 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07674 3007 4413 3006 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07673 3006 5225 3007 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07672 7514 3514 3515 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07671 3514 5000 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07670 3515 4673 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07669 7514 3820 1010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07668 1010 2591 1043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07667 1500 1043 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07666 7514 6468 6469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07665 6468 6532 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07664 6469 6954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07663 2577 2926 2579 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07662 2579 3135 2578 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07661 2578 3499 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07660 2575 2925 2579 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07659 7514 5137 2575 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07658 7514 6025 2577 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07657 2576 2579 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07656 7514 1851 1225 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07655 1225 1883 1277 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07654 1558 1277 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07653 7514 4005 4006 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07652 4005 6133 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07651 4006 6846 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07650 4023 5001 4024 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07649 4024 5718 4073 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07648 7514 5000 4023 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07647 4149 4073 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07646 7514 1759 1761 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07645 1761 2037 1760 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07644 1973 1760 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07643 7514 4695 2484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07642 2484 2590 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07641 2514 2515 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07640 2484 4697 2515 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07639 2515 2517 2484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07638 6784 6828 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07637 6782 6830 6822 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07636 7514 7481 6782 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07635 7514 7208 6830 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07634 6829 6830 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07633 7514 6825 6828 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07632 6824 6827 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07631 7514 6824 6783 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07630 6822 6829 6824 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07629 7481 6822 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07628 7514 6822 7481 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07627 6783 6829 6827 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07626 6827 6830 6784 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07625 7057 7086 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07624 7055 7088 7082 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07623 7514 7464 7055 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07622 7514 7199 7088 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07621 7089 7088 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07620 7514 7084 7086 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07619 7083 7085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07618 7514 7083 7056 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07617 7082 7089 7083 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07616 7464 7082 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07615 7514 7082 7464 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07614 7056 7089 7085 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07613 7085 7088 7057 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07612 793 1572 753 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07611 753 1046 793 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07610 7514 979 753 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07609 6027 6165 6028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07608 6028 6166 6027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07607 7514 6125 6028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07606 7358 7357 7359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07605 7359 7458 7358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07604 7514 7420 7359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07603 5334 5502 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07602 5353 5352 5334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07601 5412 5411 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07600 5500 7010 5412 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07599 2571 3023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07598 2991 2591 2571 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07597 7514 1464 737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07596 737 1598 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07595 1548 760 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07594 737 1465 760 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07593 760 1466 737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07592 2024 2263 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07591 2154 3023 2024 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07590 264 3549 246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07589 246 3545 264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07588 7514 3546 246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07587 262 264 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07586 5422 5420 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07585 5423 5421 5422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07584 6446 7033 6447 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07583 6445 6631 6446 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07582 6447 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07581 6444 6446 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07580 7514 7032 6445 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07579 6445 7129 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07578 6916 7391 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07577 6917 7384 6916 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07576 5767 6968 5768 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07575 5768 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07574 5804 7454 5767 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07573 6021 7491 6020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07572 6020 7379 6021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07571 7514 6628 6020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07570 6160 6021 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07569 5605 5981 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07568 7514 5818 5605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07567 5605 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07566 7514 5815 5605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07565 5604 5605 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07564 6531 6565 6505 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07563 6505 6566 6531 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07562 7514 7452 6505 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07561 3056 4600 3057 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07560 3057 4603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07559 3055 5841 3056 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07558 4568 6333 3055 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07557 6714 6652 6062 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07556 7514 6061 6063 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07555 6062 6063 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07554 7514 4695 2202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07553 2202 2442 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07552 2241 2242 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07551 2202 4697 2242 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07550 2242 2245 2202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07549 6940 7075 6918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07548 6918 7255 6940 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07547 7514 7420 6918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07546 3357 4158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07545 3356 3515 3357 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07544 3355 5043 3356 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07543 7514 3922 3355 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07542 3355 3925 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07541 4894 5841 4895 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07540 4895 5691 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07539 5252 5690 4894 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07538 2425 2842 2057 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07537 2057 2792 2425 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07536 7514 2504 2057 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07535 7514 1851 1853 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07534 1853 2576 1854 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07533 1852 1854 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07532 6449 6676 6448 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07531 6448 6869 6450 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07530 7514 6965 6449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07529 6553 6450 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07528 4468 4732 4469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07527 4469 5093 4510 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07526 7514 5178 4468 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07525 4585 4510 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07524 5643 5895 5642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07523 5642 5678 5680 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07522 7514 5679 5643 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07521 5677 5680 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07520 577 653 578 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07519 578 833 577 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07518 7514 778 578 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07517 576 577 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07516 2002 2009 1731 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07515 1731 2007 2002 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07514 7514 2008 1731 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07513 3258 3665 3201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07512 3201 3738 3258 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07511 7514 3513 3201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07510 3256 3258 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07509 5848 5917 5790 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07508 5790 6058 5848 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07507 7514 5846 5790 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07506 6010 7491 5865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07505 5865 7379 6010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07504 7514 7335 5865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07503 7514 3023 2201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07502 2201 2263 2236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07501 2292 2236 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07500 7456 7461 7458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07499 7514 7455 7456 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07498 7459 7460 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07497 7458 7457 7459 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07496 7514 7460 7461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07495 7457 7455 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07494 7289 7387 7288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07493 7288 7513 7289 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07492 7514 7287 7288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07491 6389 6393 6354 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07490 6354 6394 6389 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07489 7514 6388 6354 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07488 7514 1500 1133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07487 1133 1501 1164 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07486 2543 1164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07485 5935 5988 5936 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07484 5936 5989 5990 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07483 7514 6044 5935 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07482 5987 5990 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07481 7514 6408 6217 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07480 6217 6407 6260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07479 6474 6260 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07478 7514 4376 758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07477 758 3820 797 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07476 2880 797 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07475 216 1466 215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07474 215 461 216 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07473 7514 511 215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07472 507 216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07471 1518 1559 1556 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07470 7514 1560 1518 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07469 1519 1558 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07468 1556 1555 1519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07467 7514 1558 1559 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07466 1555 1560 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07465 7113 7496 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07464 5225 5138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07463 534 536 493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07462 493 533 534 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07461 7514 4600 493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07460 4728 534 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07459 4333 4447 4334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07458 4334 4448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07457 4332 5173 4333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07456 5994 4375 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07455 4375 4446 4332 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07454 3249 3420 3199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07453 3199 3917 3249 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07452 7514 4823 3199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07451 3248 3249 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07450 3361 3398 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07449 3359 3402 3394 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07448 7514 3696 3359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07447 7514 3400 3402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07446 3401 3402 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07445 7514 3695 3398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07444 3396 3397 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07443 7514 3396 3360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07442 3394 3401 3396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07441 3696 3394 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07440 7514 3394 3696 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07439 3360 3401 3397 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07438 3397 3402 3361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07437 7136 7139 7137 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07436 7514 7464 7136 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07435 7138 7418 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07434 7137 7135 7138 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07433 7514 7418 7139 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07432 7135 7464 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07431 7514 5385 5378 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07430 5378 6846 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07429 7514 5467 5378 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07428 2353 4724 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07427 2929 5889 2353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07426 7201 7491 7177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07425 7177 7379 7201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07424 7514 7462 7177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07423 7261 7201 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07422 7514 3601 3544 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07421 3544 3666 3602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07420 4172 3602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07419 2573 2684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07418 2613 2814 2573 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07417 1428 1823 1397 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07416 1397 3545 1428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07415 7514 3546 1397 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07414 1427 1428 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07413 7047 7391 7048 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07412 7048 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07411 7046 7113 7047 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07410 7045 7114 7046 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07409 5880 5966 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07408 5881 5879 5880 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07407 7514 6432 3976 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07406 3976 5128 4035 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07405 7514 5128 4033 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07404 4035 4033 3977 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07403 6439 4035 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07402 3977 4574 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07401 7514 6617 3621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07400 3621 5128 3623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07399 7514 5128 3622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07398 3623 3622 3624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07397 6620 3623 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07396 3624 3870 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07395 7514 3550 3297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07394 3297 5128 3296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07393 7514 5128 3299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07392 3296 3299 3298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07391 3554 3296 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07390 3298 4217 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07389 744 1155 745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07388 745 775 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07387 776 1688 744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07386 2302 2383 2303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07385 2303 2514 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07384 2424 2304 2302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07383 7514 5156 5157 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07382 5157 5158 5159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07381 5830 5159 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07380 1541 4377 1542 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07379 1542 1707 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07378 1540 5173 1541 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07377 1581 4376 1540 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07376 2636 5001 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07375 2739 5840 2636 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07374 2635 2816 2739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07373 7514 2679 2635 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07372 2634 5842 2739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07371 7514 7108 2634 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07370 1240 1915 1239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07369 1239 1384 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07368 1624 3742 1240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07367 6774 6849 6775 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07366 6775 7049 6774 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07365 7514 6917 6775 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07364 6773 6774 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07363 7476 7475 7478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07362 7478 7477 7479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07361 7514 7480 7476 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07360 7474 7479 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07359 4317 4979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07358 4771 5832 4317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07357 7514 4425 4771 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07356 4450 4447 4451 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07355 4451 4448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07354 4449 5173 4450 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07353 4789 4446 4449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07352 4398 4437 4399 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07351 4399 4600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07350 4397 5841 4398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07349 4995 4433 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07348 4433 6333 4397 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07347 2334 2332 2336 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07346 2336 2463 2335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07345 7514 2333 2334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07344 3033 2335 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07343 442 479 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07342 438 444 478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07341 7514 437 438 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07340 7514 669 444 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07339 443 444 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07338 7514 480 479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07337 439 440 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07336 7514 439 441 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07335 478 443 439 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07334 437 478 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07333 7514 478 437 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07332 441 443 440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07331 440 444 442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07330 561 819 560 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07329 560 765 562 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07328 7514 1809 561 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07327 696 562 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07326 7514 5275 5351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07325 5351 4715 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07324 7514 5273 5351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07323 3920 4158 3863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07322 7514 4156 3921 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07321 3863 3921 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07320 7514 1373 1041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07319 1041 975 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07318 7514 1044 1041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07317 1670 4600 1671 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07316 1671 2033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07315 1669 2103 1670 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07314 2946 1703 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07313 1703 7162 1669 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07312 2860 3501 2859 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07311 2859 4669 2860 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07310 7514 2949 2859 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07309 4610 4760 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07308 4641 4762 4610 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07307 4974 5056 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07306 4973 6444 4974 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07305 7514 6538 5626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07304 5626 5625 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07303 7514 5909 5626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07302 7514 5720 5846 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07301 5846 6538 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07300 7514 5909 5846 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07299 7375 7374 7377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07298 7514 7488 7375 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07297 7378 7486 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07296 7377 7376 7378 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07295 7514 7486 7374 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07294 7376 7488 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07293 7256 7280 7257 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07292 7257 7428 7256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07291 7514 7453 7257 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07290 7255 7256 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07289 4810 4982 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07288 5515 4809 4810 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07287 7514 3179 2879 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07286 2879 3178 2878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07285 3116 2878 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07284 6803 7168 6802 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07283 6802 6912 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07282 6851 7387 6803 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07281 7514 2608 2610 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07280 2610 2612 2609 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07279 5128 2609 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07278 5339 5364 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07277 5365 6099 5339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07276 1406 1619 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07275 2220 1620 1406 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07274 1405 1834 2220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07273 7514 3425 1405 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07272 1405 1631 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07271 7043 7042 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07270 7044 7109 7043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07269 7041 7384 7044 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07268 7514 7286 7041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07267 7041 7391 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07266 3994 4215 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07265 5681 4228 3994 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07264 3995 3993 5681 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07263 7514 4149 3995 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07262 3995 5909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07261 6798 7110 6799 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07260 6799 6843 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07259 7381 6907 6798 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07258 7514 4926 4882 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07257 4882 4927 4928 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07256 5243 4928 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07255 2836 3418 2702 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07254 2702 2929 2836 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07253 7514 6388 2702 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07252 1362 2174 1361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07251 1361 1837 1362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07250 7514 7162 1361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07249 1431 1362 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07248 2470 2880 2469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07247 2469 2684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07246 2468 4446 2470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07245 2467 2881 2468 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07244 2068 2880 2069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07243 2069 2263 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07242 2067 4446 2068 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07241 2337 2881 2067 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07240 211 214 894 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07239 7514 462 211 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07238 213 1021 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07237 894 212 213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07236 7514 1021 214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07235 212 462 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07234 5778 5833 5777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07233 5777 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07232 5776 5841 5778 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07231 6128 7162 5776 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07230 7258 7464 7260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07229 7260 7418 7259 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07228 7514 7462 7258 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07227 7460 7259 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07226 5415 5413 5414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07225 5414 7358 5416 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07224 7514 5804 5415 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07223 5505 5416 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07222 2797 3149 2761 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07221 2761 4695 2797 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07220 7514 2856 2761 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07219 2795 2797 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07218 7514 2837 2195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07217 2195 2785 2212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07216 2287 2212 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07215 7514 1851 249 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07214 249 2696 271 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07213 272 271 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07212 7514 2811 1940 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07211 1940 1971 1972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07210 1970 1972 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07209 3097 3501 3049 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07208 3049 4669 3097 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07207 7514 3499 3049 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07206 5861 5864 6014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07205 7514 5860 5861 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07204 5863 6726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07203 6014 5862 5863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07202 7514 6726 5864 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07201 5862 5860 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07200 7099 7491 7063 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07199 7063 7379 7099 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07198 7514 7489 7063 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07197 5445 5448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07196 5441 5450 5443 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07195 7514 5536 5441 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07194 7514 5449 5450 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07193 5447 5450 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07192 7514 5535 5448 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07191 5442 5444 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07190 7514 5442 5446 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07189 5443 5447 5442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07188 5536 5443 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07187 7514 5443 5536 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07186 5446 5447 5444 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07185 5444 5450 5445 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07184 4762 5884 4735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07183 4735 5885 4762 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07182 7514 5069 4735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07181 5478 5516 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07180 5476 5519 5510 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07179 7514 7511 5476 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07178 7514 5518 5519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07177 5517 5519 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07176 7514 5515 5516 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07175 5511 5513 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07174 7514 5511 5477 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07173 5510 5517 5511 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07172 7511 5510 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07171 7514 5510 7511 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07170 5477 5517 5513 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07169 5513 5519 5478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07168 2074 2800 2073 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07167 2073 2300 2089 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07166 7514 2801 2074 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07165 2088 2089 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07164 2245 2596 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07163 1284 1092 1093 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07162 1093 1091 1284 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07161 7514 1159 1093 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07160 3839 3837 3838 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07159 3838 4673 3839 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07158 7514 6576 3838 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07157 3836 3839 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07156 7014 7034 7013 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07155 7012 7078 7014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07154 7013 7033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07153 7010 7014 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07152 7514 7032 7012 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07151 7012 7011 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_07150 5171 1449 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07149 7514 1168 5171 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07148 4852 4979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07147 2590 3086 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07146 3001 6173 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07145 1885 3545 1886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07144 1886 2027 1885 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07143 7514 2029 1886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07142 3655 1885 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07141 477 528 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07140 475 530 522 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07139 7514 1449 475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07138 7514 598 530 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07137 529 530 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_07136 7514 527 528 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_07135 523 526 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07134 7514 523 476 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07133 522 529 523 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07132 1449 522 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07131 7514 522 1449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07130 476 529 526 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07129 526 530 477 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07128 254 281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07127 280 647 254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07126 253 470 280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07125 7514 468 253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07124 253 469 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07123 1871 2661 1787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07122 1787 2658 1871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07121 7514 2504 1787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07120 5817 5746 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07119 7514 2618 1114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07118 1114 1382 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07117 7514 1312 1114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07116 3142 2149 2150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07115 2150 2154 3142 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07114 7514 2164 2150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07113 1884 1883 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07112 2960 1880 1884 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07111 1882 1881 2960 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07110 7514 5735 1882 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07109 1882 5734 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07108 6734 6738 6736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07107 7514 6733 6734 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07106 6737 6819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07105 6736 6735 6737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07104 7514 6819 6738 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07103 6735 6733 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07102 7514 2541 1629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07101 1629 2543 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07100 1627 1657 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07099 1629 1628 1657 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07098 1657 2542 1629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07097 5472 5727 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07096 5797 5503 5472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07095 7514 2664 2354 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07094 2354 4106 2386 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07093 7514 4106 2387 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07092 2386 2387 2355 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07091 2669 2386 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07090 2355 3389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07089 7514 6804 3972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07088 3972 4106 3973 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07087 7514 4106 3974 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07086 3973 3974 3975 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07085 6811 3973 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07084 3975 4574 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07083 1139 1976 1138 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07082 1138 2591 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07081 1137 3820 1139 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07080 1377 4376 1137 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07079 7514 6846 4596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07078 4596 4593 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07077 4783 4595 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07076 4596 4594 4595 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07075 4595 5385 4596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_07074 1798 1833 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07073 1834 7114 1798 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07072 7514 3868 3844 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07071 3844 4106 3875 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07070 7514 4106 3871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07069 3875 3871 3845 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07068 3876 3875 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07067 3845 3870 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07066 7514 3774 3628 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07065 3628 4106 3630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07064 7514 4106 3631 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07063 3630 3631 3629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07062 3779 3630 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07061 3629 4217 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_07060 5437 7027 5440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07059 5440 5438 5439 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07058 7514 5604 5437 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07057 5670 5439 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07056 5471 6714 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07055 7514 5470 5471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07054 5471 5544 5625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07053 5625 5695 5471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07052 7172 7173 7175 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07051 7175 7174 7176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07050 7514 7287 7172 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07049 7243 7176 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07048 6382 6736 6351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07047 6351 6523 6382 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07046 7514 7420 6351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07045 1363 1365 866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07044 866 1501 1363 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07043 7514 1500 866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07042 2756 3134 2787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07041 2787 2991 2757 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07040 2757 2995 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07039 2755 2837 2787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07038 7514 2785 2755 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07037 7514 3878 2756 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07036 2784 2787 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07035 49 80 78 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07034 7514 275 49 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07033 48 771 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07032 78 77 48 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07031 7514 771 80 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07030 77 275 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_07029 7008 7464 7009 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07028 7009 7418 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07027 7007 7454 7008 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07026 7074 7015 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_07025 7015 7462 7007 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_07024 7514 3084 3045 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07023 3045 3083 3085 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07022 3636 3085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07021 1121 1342 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07020 1149 1340 1121 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07019 1120 1341 1149 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07018 7514 1551 1120 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07017 1120 1741 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_07016 7514 3412 3364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07015 3364 3411 3413 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07014 3410 3413 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07013 4617 5138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07012 5233 5832 4617 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07011 7514 4651 5233 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07010 7514 2249 2263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07009 2249 4934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07008 2263 4158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07007 1941 1973 1942 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07006 1942 1974 1975 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07005 7514 2454 1941 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07004 4360 1975 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_07003 7514 3820 1097 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07002 1097 2392 1098 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07001 1366 1098 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_07000 1807 3023 1779 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06999 1778 2292 1807 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06998 1779 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06997 3066 1807 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06996 7514 2287 1778 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06995 1778 2922 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06994 1494 1496 1495 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06993 1495 1825 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06992 1492 2315 1494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06991 1565 1493 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06990 1493 1826 1492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06989 6460 6461 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06988 6455 6463 6456 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06987 7514 7493 6455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06986 7514 6693 6463 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06985 6462 6463 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06984 7514 6466 6461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06983 6457 6458 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06982 7514 6457 6459 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06981 6456 6462 6457 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06980 7493 6456 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06979 7514 6456 7493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06978 6459 6462 6458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06977 6458 6463 6460 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06976 3383 4869 3384 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06975 3384 3432 3433 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06974 7514 3670 3383 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06973 3431 3433 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06972 2427 2431 2430 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06971 2430 2429 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06970 2428 2425 2427 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06969 3083 2426 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06968 2426 2844 2428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06967 854 896 1075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06966 7514 1809 854 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06965 855 1149 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06964 1075 897 855 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06963 7514 1149 896 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06962 897 1809 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06961 5506 5884 5190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06960 5190 5885 5506 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06959 7514 5876 5190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06958 6301 6304 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06957 6297 6305 6296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06956 7514 7475 6297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06955 7514 6302 6305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06954 6303 6305 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06953 7514 6594 6304 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06952 6298 6300 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06951 7514 6298 6299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06950 6296 6303 6298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06949 7475 6296 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06948 7514 6296 7475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06947 6299 6303 6300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06946 6300 6305 6301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06945 4671 4828 4623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06944 4622 7162 4671 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06943 4623 6266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06942 4669 4671 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06941 7514 4790 4622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06940 4622 5016 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06939 7514 4759 4760 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06938 4759 4978 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06937 4760 4973 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06936 4425 4424 4426 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06935 4426 5381 4425 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06934 7514 6386 4426 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06933 1006 1041 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06932 1091 1040 1006 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06931 7156 7227 7157 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06930 7157 7228 7156 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06929 7514 7481 7157 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06928 1560 1823 1520 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06927 1520 3545 1560 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06926 7514 3546 1520 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06925 5036 6407 5035 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06924 5035 5837 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06923 5092 6408 5036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06922 6921 6968 6920 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06921 6920 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06920 6947 7464 6921 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06919 884 1577 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06918 1371 4158 884 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06917 6408 1579 1539 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06916 1539 1765 6408 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06915 7514 1906 1539 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06914 1723 1892 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06913 7514 1753 1723 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06912 1723 2945 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06911 7514 2946 1723 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06910 2874 2958 2873 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06909 2873 2988 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06908 4824 2956 2874 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06907 836 4588 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06906 1092 4589 836 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06905 1675 4597 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06904 1764 1709 1675 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06903 2861 2945 2768 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06902 2768 2946 2861 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06901 7514 5043 2768 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06900 1788 3135 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06899 1869 3012 1788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06898 5348 5695 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06897 7514 5544 5348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06896 5348 5466 5720 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06895 5720 5467 5348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06894 6037 6393 6036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06893 6036 6394 6037 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06892 7514 6035 6036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06891 565 568 567 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06890 567 566 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06889 564 563 565 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06888 2731 2954 2732 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06887 2732 2730 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06886 2729 2743 2731 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06885 4577 2728 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06884 2728 2727 2729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06883 2022 2949 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06882 2023 3135 2022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06881 2021 2926 2023 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06880 7514 5882 2021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06879 2020 2925 2023 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06878 7514 5138 2020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06877 5343 5891 5344 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06876 5344 5992 5370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06875 7514 5889 5343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06874 5369 5370 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06873 5638 5662 5639 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06872 5639 7263 5663 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06871 7514 6023 5638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06870 5809 5663 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06869 1077 1074 1076 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06868 1076 1075 1078 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06867 7514 1145 1077 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06866 1267 1078 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06865 7029 7033 7030 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06864 7028 7099 7029 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06863 7030 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06862 7027 7029 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06861 7514 7032 7028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06860 7028 7484 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06859 7514 6897 6359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06858 6359 6400 6398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06857 6397 6398 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06856 7514 3632 3635 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06855 3635 3633 3634 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06854 4265 3634 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06853 7514 3240 1649 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06852 1744 1649 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06851 7514 1649 1744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06850 7514 1649 1744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06849 1744 1649 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06848 7514 1744 1278 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06847 3081 1278 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06846 7514 1278 3081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06845 7514 1278 3081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06844 3081 1278 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06843 7514 1744 1745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06842 3135 1745 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06841 7514 1745 3135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06840 7514 1745 3135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06839 3135 1745 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06838 7514 286 287 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06837 390 287 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06836 7514 287 390 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06835 7514 287 390 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06834 390 287 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06833 7514 390 189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06832 2686 189 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06831 7514 189 2686 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06830 7514 189 2686 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06829 2686 189 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06828 7514 390 391 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06827 4158 391 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06826 7514 391 4158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06825 7514 391 4158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06824 4158 391 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06823 644 823 621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06822 621 824 644 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06821 7514 900 621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06820 698 644 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06819 1616 1652 1615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06818 1615 1653 1651 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06817 7514 1828 1616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06816 4695 1651 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06815 1012 1047 1013 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06814 1013 1376 1048 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06813 7514 1363 1012 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06812 1046 1048 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06811 7514 1449 608 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06810 608 1168 607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06809 1052 607 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06808 5211 5454 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06807 3978 6025 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06806 3770 6804 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06805 4423 5889 4422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06804 4421 4986 4423 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06803 4422 4589 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06802 6246 4423 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06801 7514 4987 4421 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06800 4421 4984 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06799 277 280 252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06798 252 276 277 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06797 7514 512 252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06796 899 277 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06795 4908 5216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06794 4698 5125 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06793 4121 4120 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06792 4114 4122 4115 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06791 7514 4113 4114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06790 7514 4488 4122 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06789 4123 4122 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06788 7514 4119 4120 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06787 4116 4118 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06786 7514 4116 4117 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06785 4115 4123 4116 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06784 4113 4115 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06783 7514 4115 4113 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06782 4117 4123 4118 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06781 4118 4122 4121 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06780 3259 3922 3202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06779 3202 3925 3259 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06778 7514 5216 3202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06777 2454 2543 2065 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06776 2065 2541 2454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06775 7514 2322 2065 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06774 1802 4000 1803 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06773 1803 1837 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06772 2182 6333 1802 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06771 7183 7286 7184 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06770 7184 7356 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06769 7234 7384 7183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06768 5664 6029 5631 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06767 5631 6030 5664 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06766 7514 6125 5631 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06765 7514 4424 3325 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06764 3325 4264 3327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06763 7514 4264 3329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06762 3327 3329 3328 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06761 3324 3327 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06760 3328 3326 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06759 7514 4718 3807 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06758 3807 4264 3806 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06757 7514 4264 3809 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06756 3806 3809 3808 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06755 3905 3806 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06754 3808 6894 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06753 7514 4991 3195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06752 3195 4264 3224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06751 7514 4264 3225 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06750 3224 3225 3194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06749 3568 3224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06748 3194 3300 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06747 6789 6836 6790 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06746 6790 7098 6838 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06745 7514 6837 6789 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06744 6892 6838 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06743 6664 6698 6665 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06742 6665 7149 6699 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06741 7514 6696 6664 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06740 6697 6699 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06739 1648 2101 1647 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06738 1647 2241 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06737 1699 2165 1648 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06736 7514 4431 3677 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06735 3677 4264 3712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06734 7514 4264 3715 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06733 3712 3715 3678 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06732 3953 3712 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06731 3678 3713 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_06730 859 3814 858 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06729 858 2174 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06728 857 4158 859 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06727 1809 5690 857 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06726 3381 5173 3380 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06725 3380 5172 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06724 3379 4446 3381 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06723 4673 3742 3379 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06722 5284 5282 5283 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06721 5283 6015 5285 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06720 7514 6017 5284 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06719 5507 5285 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06718 7514 2662 2629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06717 2629 3156 2663 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06716 3128 2663 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06715 7514 2602 1903 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06714 1903 2536 1902 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06713 2039 1902 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06712 1478 1851 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06711 1479 1876 1478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06710 1477 1688 1479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06709 7514 2095 1477 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06708 1477 3545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06707 1861 2007 1862 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06706 1862 1860 1861 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06705 7514 2009 1862 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06704 4984 1861 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06703 7052 7077 7075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06702 7514 7196 7052 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06701 7053 7074 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06700 7075 7073 7053 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06699 7514 7074 7077 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06698 7073 7196 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06697 7514 1271 1223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06696 1223 1809 1272 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06695 1270 1272 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06694 7514 6980 3171 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06693 3171 6979 3172 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06692 3170 3172 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06691 7514 2948 2858 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06690 2858 3232 2857 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06689 2856 2857 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06688 710 778 712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06687 712 777 711 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06686 7514 776 710 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06685 709 711 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06684 515 468 432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06683 432 469 515 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06682 7514 470 432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06681 1773 4600 1772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06680 1772 4603 1774 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06679 7514 6133 1773 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06678 1771 1774 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06677 2311 2313 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06676 2306 2314 2307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06675 7514 2596 2306 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06674 7514 2672 2314 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06673 2312 2314 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06672 7514 2597 2313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06671 2308 2309 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06670 7514 2308 2310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06669 2307 2312 2308 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06668 2596 2307 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06667 7514 2307 2596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06666 2310 2312 2309 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06665 2309 2314 2311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06664 1212 1915 1213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06663 1213 1384 1241 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06662 7514 3742 1212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06661 1211 1241 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06660 6786 6968 6785 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06659 6785 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06658 6831 7466 6786 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06657 3729 5541 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06656 7514 3456 3729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06655 3729 5377 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06654 7514 5378 3729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06653 4651 4504 4462 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06652 4462 5381 4651 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06651 7514 6386 4462 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06650 1507 4597 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06649 1765 1624 1507 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06648 7514 7390 6854 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06647 6854 7388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06646 6852 6854 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06645 6052 6112 6053 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06644 6053 6336 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06643 6393 6576 6052 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06642 6315 5617 5618 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06641 5618 5616 6315 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06640 7514 5889 5618 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06639 1467 1464 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06638 7514 1598 1467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06637 1467 1465 1810 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06636 1810 1466 1467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06635 1399 1430 1400 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06634 1400 1723 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06633 1881 1466 1399 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06632 7514 7453 6495 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06631 6495 7074 6550 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06630 6518 6550 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06629 7514 4365 4912 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06628 4365 4364 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06627 4912 6600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06626 2778 6339 2777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06625 2777 4296 2821 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06624 7514 2820 2778 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06623 2819 2821 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06622 6201 6202 6204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06621 6204 7242 6203 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06620 7514 7111 6201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06619 6272 6203 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06618 2011 2009 2010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06617 2010 2007 2011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06616 7514 2008 2010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06615 2081 2011 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06614 5927 5967 5926 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06613 5926 6382 5968 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06612 7514 6102 5927 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06611 5966 5968 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06610 7514 3958 3639 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06609 7514 3957 3639 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06608 3639 6030 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06607 4211 3639 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06606 5920 5949 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06605 5918 5951 5944 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06604 7514 7453 5918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06603 7514 6231 5951 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06602 5950 5951 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06601 7514 5954 5949 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06600 5945 5948 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06599 7514 5945 5919 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06598 5944 5950 5945 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06597 7453 5944 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06596 7514 5944 7453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06595 5919 5950 5948 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06594 5948 5951 5920 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06593 7514 1851 622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06592 622 2371 646 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06591 771 646 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06590 7514 6840 6645 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06589 6645 6644 6647 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06588 6646 6647 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06587 7514 1830 1797 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06586 1797 2041 1831 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06585 1832 1831 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06584 7514 4773 1795 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06583 1795 2102 1829 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06582 1828 1829 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06581 6903 7320 6905 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06580 6905 6902 6904 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06579 7514 7039 6903 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06578 6901 6904 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06577 5593 5596 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06576 5588 5597 5589 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06575 7514 6676 5588 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06574 7514 5594 5597 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06573 5595 5597 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06572 7514 5881 5596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06571 5590 5591 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06570 7514 5590 5592 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06569 5589 5595 5590 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06568 6676 5589 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06567 7514 5589 6676 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06566 5592 5595 5591 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06565 5591 5597 5593 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06564 3009 2945 2767 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06563 2767 2946 3009 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06562 7514 5274 2767 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06561 5021 5052 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06560 5019 5054 5046 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06559 7514 5045 5019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06558 7514 5270 5054 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06557 5053 5054 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06556 7514 5051 5052 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06555 5047 5050 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06554 7514 5047 5020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06553 5046 5053 5047 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06552 5045 5046 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06551 7514 5046 5045 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06550 5020 5053 5050 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06549 5050 5054 5021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06548 1794 2315 1793 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06547 1793 1825 1827 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06546 7514 1826 1794 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06545 2288 1827 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06544 7514 1915 1214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06543 1214 1908 1242 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06542 1579 1242 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06541 4197 6388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06540 5547 5553 5548 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06539 5494 5555 5547 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06538 6061 5547 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06537 7514 5547 6061 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06536 5497 5552 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06535 7514 5848 5552 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06534 5553 5555 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06533 7514 5554 5555 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06532 5495 5550 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06531 5548 7500 5495 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06530 5550 5555 5497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06529 5496 5553 5550 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06528 7514 5548 5496 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06527 7514 6061 5493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06526 5493 7500 5494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06525 5606 5523 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06524 3705 5887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06523 5981 6187 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06522 7514 6040 6041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06521 6040 6039 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06520 6041 6111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06519 2072 2120 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06518 2070 2121 2113 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06517 7514 2111 2070 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06516 7514 2553 2121 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06515 2119 2121 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06514 7514 2118 2120 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06513 2114 2117 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06512 7514 2114 2071 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06511 2113 2119 2114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06510 2111 2113 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06509 7514 2113 2111 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06508 2071 2119 2117 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06507 2117 2121 2072 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06506 3830 3663 3664 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06505 3664 6340 3830 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06504 7514 3737 3664 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06503 634 4934 635 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06502 635 3820 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06501 633 1449 634 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06500 1908 672 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06499 672 4376 633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06498 4255 6392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06497 5051 6894 4402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06496 4402 4401 5051 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06495 7514 4629 4402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06494 4883 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06493 5226 7286 4883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06492 7212 7210 7179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06491 7179 7270 7212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06490 7514 7420 7179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06489 7514 6386 6320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06488 6320 6318 6319 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06487 6836 6319 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06486 3957 2088 2019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06485 2019 2153 3957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06484 7514 2018 2019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06483 6514 6912 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06482 6534 7168 6514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06481 7514 5082 5034 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06480 5034 5083 5084 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06479 5678 5084 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06478 7433 7334 7282 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06477 7282 7383 7433 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06476 7514 7453 7282 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06475 4184 4427 4185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06474 4185 4231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06473 4183 4370 4184 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06472 4364 4225 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06471 4225 4224 4183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06470 7514 7285 7286 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06469 7285 7390 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06468 7286 7388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06467 1932 2241 1933 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06466 1933 2023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06465 1931 2101 1932 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06464 1967 2165 1931 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06463 3658 4588 3661 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06462 3661 3660 3662 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06461 7514 4724 3658 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06460 3659 3662 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06459 512 3081 487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06458 487 1187 512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06457 7514 906 487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06456 3075 3074 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06455 7514 3069 3075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06454 3075 3070 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06453 7514 3071 3075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06452 6169 3075 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06451 7514 6344 2356 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06450 2356 2743 2388 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06449 2676 2388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06448 7514 2653 2624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06447 2624 2652 2654 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06446 2655 2654 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06445 2346 2926 2373 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06444 2373 3081 2347 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06443 2347 3226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06442 2345 2925 2373 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06441 7514 5274 2345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06440 7514 5887 2346 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06439 2371 2373 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06438 1962 2792 1924 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06437 1924 2842 1962 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06436 7514 2371 1924 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06435 2149 1962 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06434 6358 6914 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06433 6698 6529 6358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06432 6357 6392 6698 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06431 7514 6393 6357 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06430 6357 6394 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06429 1100 3820 1099 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06428 1099 2591 1101 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06427 7514 2881 1100 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06426 1368 1101 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06425 1632 1838 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06424 7514 1771 1632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06423 4314 4353 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06422 4312 4355 4347 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06421 7514 5882 4312 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06420 7514 4488 4355 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06419 4354 4355 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06418 7514 4416 4353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_06417 4350 4352 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06416 7514 4350 4313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06415 4347 4354 4350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06414 5882 4347 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06413 7514 4347 5882 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06412 4313 4354 4352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06411 4352 4355 4314 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06410 962 1700 961 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06409 961 1968 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06408 959 1435 962 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06407 960 958 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06406 958 4368 959 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06405 1004 1700 1003 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06404 1003 1968 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06403 1002 1435 1004 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06402 1037 1038 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06401 1038 1688 1002 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06400 1577 1709 1538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06399 1538 1624 1577 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06398 7514 4597 1538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06397 3970 4448 3971 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06396 3971 4441 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06395 3969 4442 3970 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06394 5691 4004 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06393 4004 4934 3969 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06392 4740 5055 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06391 5158 5832 4740 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06390 7514 4862 5158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06389 6964 7280 6919 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06388 6919 7428 6964 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06387 7514 6965 6919 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06386 6942 6964 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06385 6883 6968 6881 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06384 6881 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06383 6882 7475 6883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06382 6151 7034 6153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06381 6152 6519 6151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06380 6153 7033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06379 6150 6151 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06378 7514 7032 6152 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06377 6152 6291 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06376 221 224 907 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06375 7514 225 221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06374 223 576 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06373 907 222 223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06372 7514 576 224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06371 222 225 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06370 2291 3135 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06369 2290 3499 2291 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06368 4896 6135 4897 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06367 4897 4938 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06366 7242 4937 4896 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06365 7514 6839 6213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06364 6213 6648 6252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06363 6386 6252 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06362 6896 6980 6898 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06361 6898 6979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06360 6897 7481 6896 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06359 2304 3418 2305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06358 2305 2929 2304 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06357 7514 6173 2305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06356 1563 3023 1522 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06355 1521 2292 1563 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06354 1522 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06353 1965 1563 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06352 7514 2159 1521 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06351 1521 2095 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_06350 7514 2820 2749 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06349 2749 6339 2750 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06348 2751 2750 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06347 7514 2708 649 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06346 649 1037 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06345 647 649 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06344 7514 974 2591 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06343 974 2686 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06342 2591 4934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06341 7514 6333 3518 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06340 3518 5623 3517 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06339 3516 3517 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06338 6519 7491 6496 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06337 6496 7379 6519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06336 7514 7452 6496 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06335 7514 3957 3983 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06334 3983 3958 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06333 6029 3983 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06332 1370 4437 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06331 1369 1368 1370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06330 1367 1365 1369 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06329 7514 1366 1367 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06328 1367 1500 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06327 7514 5378 3243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06326 7514 5541 3243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06325 3243 5377 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06324 3240 3243 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06323 24 25 370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06322 7514 78 24 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06321 26 126 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06320 370 23 26 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06319 7514 126 25 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06318 23 78 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06317 3349 3347 3350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06316 3350 4372 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06315 3345 3348 3349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06314 3346 3344 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_06313 3344 3343 3345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06312 3311 3319 3312 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06311 3308 3318 3311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06310 4502 3311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06309 7514 3311 4502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06308 3316 3317 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06307 7514 3315 3317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06306 3319 3318 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06305 7514 3571 3318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06304 3310 3314 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06303 3312 5100 3310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06302 3314 3318 3316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06301 3313 3319 3314 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06300 7514 3312 3313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06299 7514 4502 3309 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06298 3309 5100 3308 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06297 3865 6133 3864 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06296 3864 5994 3923 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06295 7514 5000 3865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06294 3922 3923 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06293 902 3081 485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06292 485 2134 902 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06291 7514 509 485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06290 751 2816 752 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06289 752 790 791 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06288 7514 3023 751 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06287 975 791 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06286 1601 1810 1602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06285 1602 1954 1639 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06284 7514 1809 1601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06283 1860 1639 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06282 1482 2424 1483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06281 1483 1699 1484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06280 1484 2504 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06279 1481 2789 1483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06278 7514 2416 1481 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06277 7514 2502 1482 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06276 2090 1483 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06275 7514 7381 7382 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06274 7490 7382 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06273 7514 7382 7490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06272 7514 7382 7490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06271 7490 7382 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06270 7514 7490 7281 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06269 7280 7281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06268 7514 7281 7280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06267 7514 7281 7280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06266 7280 7281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06265 7514 7490 7492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06264 7491 7492 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06263 7514 7492 7491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06262 7514 7492 7491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06261 7491 7492 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06260 6658 6876 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06259 7084 6681 6658 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06258 831 2300 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06257 7514 1037 831 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06256 632 3352 631 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06255 631 3820 671 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06254 7514 4376 632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06253 1049 671 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06252 3913 3997 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06251 3710 4113 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06250 4916 5043 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06249 5543 7388 5491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06248 5491 7390 5543 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06247 7514 7384 5491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06246 5541 5543 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06245 2383 2381 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06244 7514 2810 2383 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_06243 5784 5842 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06242 5902 7108 5784 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06241 5783 5840 5902 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06240 7514 5841 5783 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06239 5783 6133 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_06238 7514 1264 311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06237 310 311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06236 7514 311 310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06235 7514 311 310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06234 310 311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06233 7514 1264 359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06232 358 359 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06231 7514 359 358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06230 7514 359 358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06229 358 359 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06228 7514 1264 361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06227 360 361 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06226 7514 361 360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06225 7514 361 360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06224 360 361 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06223 7514 1264 317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06222 316 317 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06221 7514 317 316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06220 7514 317 316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06219 316 317 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06218 7514 1264 367 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06217 366 367 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06216 7514 367 366 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06215 7514 367 366 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06214 366 367 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06213 7514 1264 369 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06212 368 369 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06211 7514 369 368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06210 7514 369 368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06209 368 369 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06208 7514 1264 1219 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06207 1180 1219 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06206 7514 1219 1180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06205 7514 1219 1180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06204 1180 1219 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06203 7424 7466 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06202 6629 6628 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06201 6195 5912 5624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06200 5624 5623 6195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06199 7514 6333 5624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06198 7514 6599 7032 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06197 7032 6848 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06196 7514 6600 7032 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06195 2791 2792 2758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06194 2758 2842 2791 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06193 7514 2789 2758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06192 3069 2791 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06191 7169 7236 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06190 7168 7287 7169 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06189 7514 1264 1254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06188 1253 1254 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06187 7514 1254 1253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06186 7514 1254 1253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06185 1253 1254 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06184 7514 1264 1256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06183 1255 1256 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06182 7514 1256 1255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06181 7514 1256 1255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06180 1255 1256 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06179 7514 1264 1222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06178 1185 1222 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06177 7514 1222 1185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06176 7514 1222 1185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06175 1185 1222 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06174 7514 1264 1262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06173 1261 1262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06172 7514 1262 1261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06171 7514 1262 1261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06170 1261 1262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06169 7514 1264 1265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06168 1263 1265 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06167 7514 1265 1263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06166 7514 1265 1263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06165 1263 1265 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06164 7514 1281 321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06163 320 321 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06162 7514 321 320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06161 7514 321 320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06160 320 321 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06159 7514 1281 375 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06158 374 375 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06157 7514 375 374 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06156 7514 375 374 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06155 374 375 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06154 7514 1281 377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06153 376 377 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06152 7514 377 376 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06151 7514 377 376 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06150 376 377 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06149 5006 5013 5008 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06148 5005 5015 5006 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06147 7235 5006 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06146 7514 5006 7235 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06145 5011 5014 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06144 7514 5012 5014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06143 5013 5015 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06142 7514 5554 5015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06141 5007 5010 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06140 5008 7500 5007 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06139 5010 5015 5011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06138 5009 5013 5010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06137 7514 5008 5009 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06136 7514 7235 5004 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06135 5004 7500 5005 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_06134 486 827 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06133 511 564 486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06132 1758 4158 1757 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06131 1757 1837 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06130 1830 7114 1758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06129 1095 2255 1096 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06128 1096 1363 1095 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06127 7514 1449 1096 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06126 1203 1095 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06125 3671 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06124 3670 5001 3671 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06123 5650 6652 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06122 5695 6061 5650 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06121 7514 6965 6781 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06120 6781 6869 6820 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06119 6819 6820 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06118 3016 3160 3015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06117 3015 3303 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06116 3017 3159 3016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06115 6340 3326 3017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06114 7514 6271 6221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06113 6221 6272 6273 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06112 6341 6273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06111 7514 7464 7360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06110 7360 7418 7361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06109 7413 7361 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06108 7514 1281 327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06107 326 327 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06106 7514 327 326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06105 7514 327 326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06104 326 327 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06103 7514 1281 383 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06102 382 383 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06101 7514 383 382 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06100 7514 383 382 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06099 382 383 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06098 7514 1281 385 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06097 384 385 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06096 7514 385 384 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06095 7514 385 384 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06094 384 385 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06093 7514 1281 1224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06092 1190 1224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06091 7514 1224 1190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06090 7514 1224 1190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06089 1190 1224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06088 7514 1281 1274 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06087 1273 1274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06086 7514 1274 1273 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06085 7514 1274 1273 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06084 1273 1274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06083 7514 1281 1276 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06082 1275 1276 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06081 7514 1276 1275 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06080 7514 1276 1275 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06079 1275 1276 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06078 7514 1281 1227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06077 1196 1227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06076 7514 1227 1196 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06075 7514 1227 1196 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06074 1196 1227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06073 7514 5752 5733 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06072 6739 5733 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06071 7514 5733 6739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06070 7514 5733 6739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06069 6739 5733 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06068 7514 5752 5753 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06067 6771 5753 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06066 7514 5753 6771 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06065 7514 5753 6771 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06064 6771 5753 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06063 7514 3717 3718 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06062 5752 3718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06061 7514 3718 5752 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06060 7514 3718 5752 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06059 5752 3718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06058 990 1025 989 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06057 989 1020 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06056 3470 1341 990 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06055 1179 1634 1178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06054 1178 1216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06053 1257 1341 1179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06052 7514 3248 2616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06051 2616 2819 2617 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06050 2884 2617 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06049 5774 7031 5775 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06048 5775 5830 5831 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06047 7514 5828 5774 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06046 5829 5831 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06045 7514 1412 736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06044 735 736 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06043 7514 736 735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06042 7514 736 735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06041 735 736 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06040 7514 735 673 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06039 5100 673 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06038 7514 673 5100 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06037 7514 673 5100 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06036 5100 673 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06035 7514 735 299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06034 7500 299 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06033 7514 299 7500 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06032 7514 299 7500 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06031 7500 299 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06030 2016 2658 2017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06029 2017 2661 2016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06028 7514 2133 2017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_06027 4280 4569 4279 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06026 4279 4568 4281 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06025 7514 4773 4280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06024 4427 4281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_06023 7514 1281 1280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06022 1279 1280 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06021 7514 1280 1279 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06020 7514 1280 1279 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06019 1279 1280 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06018 7514 1281 1283 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06017 1282 1283 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06016 7514 1283 1282 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06015 7514 1283 1282 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06014 1282 1283 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06013 7514 3210 2138 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06012 2137 2138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06011 7514 2138 2137 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06010 7514 2138 2137 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06009 2137 2138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06008 7514 3210 2214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06007 2213 2214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06006 7514 2214 2213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06005 7514 2214 2213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06004 2213 2214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06003 7514 3210 2216 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06002 2215 2216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06001 7514 2216 2215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_06000 7514 2216 2215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05999 2215 2216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05998 7514 3210 2146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05997 2145 2146 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05996 7514 2146 2145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05995 7514 2146 2145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05994 2145 2146 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05993 7514 3210 2225 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05992 2224 2225 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05991 7514 2225 2224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05990 7514 2225 2224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05989 2224 2225 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05988 7514 3210 2227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05987 2226 2227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05986 7514 2227 2226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05985 7514 2227 2226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05984 2226 2227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05983 7350 7466 7352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05982 7352 7477 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05981 7351 7475 7350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05980 7418 7367 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05979 7367 7480 7351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05978 7514 1145 994 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05977 994 1029 1030 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05976 1034 1030 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05975 3338 3663 2904 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05974 2904 2960 3338 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05973 7514 3256 2904 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05972 5200 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05971 5218 7286 5200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05970 5199 5216 5218 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05969 7514 5275 5199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05968 5199 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05967 7514 2589 2438 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05966 2438 2862 2439 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05965 2801 2439 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05964 7514 4377 4026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05963 4026 4157 4078 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05962 4077 4078 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05961 3471 3469 3473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05960 3473 3472 3474 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05959 7514 3470 3471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05958 6894 3474 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05957 3522 3559 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05956 3520 3561 3552 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05955 7514 3550 3520 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05954 7514 3558 3561 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05953 3560 3561 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05952 7514 3554 3559 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05951 3553 3556 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05950 7514 3553 3521 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05949 3552 3560 3553 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05948 3550 3552 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05947 7514 3552 3550 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05946 3521 3560 3556 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05945 3556 3561 3522 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05944 7514 2881 977 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05943 977 1384 976 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05942 1365 976 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05941 769 768 741 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05940 741 903 769 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05939 7514 1732 741 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05938 767 769 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05937 7403 7433 7402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05936 7402 7432 7434 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05935 7514 7430 7403 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05934 7431 7434 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05933 7514 2039 2041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05932 2041 2040 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05931 7514 2456 2041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05930 2638 2880 2639 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05929 2639 2684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05928 2637 4446 2638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05927 2679 2680 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05926 2680 2881 2637 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05925 6438 6440 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05924 6433 6442 6434 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05923 7514 6432 6433 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05922 7514 6622 6442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05921 6441 6442 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05920 7514 6439 6440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05919 6435 6436 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05918 7514 6435 6437 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05917 6434 6441 6435 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05916 6432 6434 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05915 7514 6434 6432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05914 6437 6441 6436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05913 6436 6442 6438 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05912 6013 7034 6012 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05911 6011 6010 6013 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05910 6012 7033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05909 6009 6013 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05908 7514 7032 6011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05907 6011 6226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05906 5640 5670 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05905 5741 5671 5640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05904 2499 2540 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05903 2738 2684 2499 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05902 1784 3646 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05901 2141 3081 1784 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05900 1783 2926 2141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05899 7514 6175 1783 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05898 1782 2925 2141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05897 7514 4834 1782 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05896 1470 1472 2082 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05895 7514 1468 1470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05894 1471 1733 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05893 2082 1469 1471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05892 7514 1733 1472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05891 1469 1468 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05890 7514 3264 3188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05889 3187 3188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05888 7514 3188 3187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05887 7514 3188 3187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05886 3187 3188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05885 7514 3264 3262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05884 3261 3262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05883 7514 3262 3261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05882 7514 3262 3261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05881 3261 3262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05880 7514 3264 3265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05879 3263 3265 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05878 7514 3265 3263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05877 7514 3265 3263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05876 3263 3265 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05875 7514 2746 865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05874 1295 865 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05873 7514 865 1295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05872 7514 865 1295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05871 1295 865 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05870 161 3346 160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05869 160 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05868 193 5841 161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05867 2890 3346 2888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05866 2888 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05865 2889 7108 2890 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05864 6874 7280 6875 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05863 6875 7428 6874 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05862 7514 7454 6875 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05861 7357 6874 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05860 6742 6968 6743 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05859 6743 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05858 6741 7481 6742 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05857 1124 1430 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05856 2133 1466 1124 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05855 765 699 620 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05854 620 698 765 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05853 7514 1341 620 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05852 1398 3135 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05851 1740 2949 1398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05850 2097 2945 2059 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05849 2059 2946 2097 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05848 7514 4979 2059 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05847 2381 2097 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05846 163 3346 164 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05845 164 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05844 162 6266 163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05843 337 3346 339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05842 339 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05841 338 6133 337 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05840 7514 2746 874 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05839 1310 874 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05838 7514 874 1310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05837 7514 874 1310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05836 1310 874 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05835 7514 2746 2726 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05834 3246 2726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05833 7514 2726 3246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05832 7514 2726 3246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05831 3246 2726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05830 7514 2746 2747 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05829 3264 2747 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05828 7514 2747 3264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05827 7514 2747 3264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05826 3264 2747 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05825 1015 4442 1016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05824 1016 1051 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05823 1111 2880 1015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05822 724 4600 723 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05821 723 1292 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05820 875 6133 724 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05819 2431 2435 2432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05818 2432 2853 2431 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05817 7514 2789 2432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05816 6335 7108 6334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05815 6334 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05814 6336 6333 6335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05813 5655 6168 5410 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05812 5410 6169 5655 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05811 7514 5876 5410 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05810 7514 5280 4194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05809 4193 4194 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05808 7514 4194 4193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05807 7514 4194 4193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05806 4193 4194 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05805 7514 5280 4246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05804 4245 4246 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05803 7514 4246 4245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05802 7514 4246 4245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05801 4245 4246 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05800 7514 5280 4248 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05799 4247 4248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05798 7514 4248 4247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05797 7514 4248 4247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05796 4247 4248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05795 7514 5280 4199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05794 4198 4199 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05793 7514 4199 4198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05792 7514 4199 4198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05791 4198 4199 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05790 7514 5280 4252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05789 4251 4252 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05788 7514 4252 4251 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05787 7514 4252 4251 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05786 4251 4252 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05785 7514 5280 4253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05784 4638 4253 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05783 7514 4253 4638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05782 7514 4253 4638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05781 4638 4253 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05780 7514 5280 5213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05779 5212 5213 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05778 7514 5213 5212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05777 7514 5213 5212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05776 5212 5213 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05775 5202 6888 5203 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05774 5203 5243 5244 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05773 7514 5241 5202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05772 5242 5244 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05771 6794 6980 6795 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05770 6795 6979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05769 6840 7489 6794 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05768 2436 2435 2437 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05767 2437 2853 2436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05766 7514 2433 2437 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05765 2434 2436 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05764 4862 4861 4863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05763 4863 5381 4862 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05762 7514 6839 4863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05761 7514 3159 3162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05760 3162 3160 3161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05759 3387 3161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05758 7514 190 192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05757 191 192 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05756 7514 192 191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05755 7514 192 191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05754 191 192 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05753 7514 191 31 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05752 7042 31 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05751 7514 31 7042 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05750 7514 31 7042 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05749 7042 31 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05748 7514 191 159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05747 5841 159 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05746 7514 159 5841 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05745 7514 159 5841 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05744 5841 159 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05743 7514 5280 5269 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05742 5268 5269 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05741 7514 5269 5268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05740 7514 5269 5268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05739 5268 5269 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05738 7514 5280 5271 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05737 5270 5271 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05736 7514 5271 5270 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05735 7514 5271 5270 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05734 5270 5271 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05733 7514 5280 5221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05732 5220 5221 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05731 7514 5221 5220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05730 7514 5221 5220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05729 5220 5221 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05728 7514 5280 5279 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05727 5278 5279 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05726 7514 5279 5278 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05725 7514 5279 5278 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05724 5278 5279 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05723 7514 5280 5281 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05722 5584 5281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05721 7514 5281 5584 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05720 7514 5281 5584 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05719 5584 5281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05718 7514 5296 4205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05717 4204 4205 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05716 7514 4205 4204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05715 7514 4205 4204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05714 4204 4205 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05713 7514 5296 4259 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05712 4258 4259 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05711 7514 4259 4258 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05710 7514 4259 4258 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05709 4258 4259 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05708 7514 5296 4260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05707 4488 4260 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05706 7514 4260 4488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05705 7514 4260 4488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05704 4488 4260 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05703 3791 3799 3792 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05702 3790 3800 3791 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05701 4861 3791 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05700 7514 3791 4861 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05699 3796 3798 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05698 7514 3797 3798 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05697 3799 3800 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05696 7514 4561 3800 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05695 3793 3795 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05694 3792 7500 3793 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05693 3795 3800 3796 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05692 3794 3799 3795 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05691 7514 3792 3794 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05690 7514 4861 3789 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05689 3789 7500 3790 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05688 6614 6344 6345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05687 6345 6410 6614 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05686 7514 6491 6345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05685 7514 4518 4471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05684 4471 4593 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05683 4517 4519 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05682 4471 4602 4519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05681 4519 5385 4471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_05680 7514 2754 1982 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05679 1981 1982 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05678 7514 1982 1981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05677 7514 1982 1981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05676 1981 1982 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05675 7514 1981 1388 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05674 5690 1388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05673 7514 1388 5690 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05672 7514 1388 5690 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05671 5690 1388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05670 7514 1981 1710 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05669 7162 1710 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05668 7514 1710 7162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05667 7514 1710 7162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05666 7162 1710 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05665 7514 1981 1582 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05664 6333 1582 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05663 7514 1582 6333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05662 7514 1582 6333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05661 6333 1582 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05660 7514 1981 1451 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05659 7114 1451 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05658 7514 1451 7114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05657 7514 1451 7114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05656 7114 1451 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05655 5924 5961 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05654 5922 5963 5955 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05653 7514 7462 5922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05652 7514 6302 5963 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05651 5964 5963 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05650 7514 5960 5961 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05649 5957 5958 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05648 7514 5957 5923 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05647 5955 5964 5957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05646 7462 5955 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05645 7514 5955 7462 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05644 5923 5964 5958 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05643 5958 5963 5924 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05642 3723 3724 3682 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05641 3682 4360 3723 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05640 7514 6397 3682 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05639 3722 3723 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05638 7514 2958 2320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05637 2320 2319 2321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05636 2318 2321 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05635 2853 3710 2852 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05634 2852 4695 2853 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05633 7514 3145 2852 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05632 7514 1449 1411 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05631 1411 4158 1450 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05630 1707 1450 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05629 7514 5296 4214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05628 4213 4214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05627 7514 4214 4213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05626 7514 4214 4213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05625 4213 4214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05624 7514 5296 4269 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05623 4268 4269 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05622 7514 4269 4268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05621 7514 4269 4268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05620 4268 4269 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05619 7514 5296 4270 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05618 4561 4270 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05617 7514 4270 4561 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05616 7514 4270 4561 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05615 4561 4270 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05614 7514 5296 5224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05613 5223 5224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05612 7514 5224 5223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05611 7514 5224 5223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05610 5223 5224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05609 7514 5296 5289 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05608 5288 5289 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05607 7514 5289 5288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05606 7514 5289 5288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05605 5288 5289 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05604 7514 5296 5290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05603 5594 5290 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05602 7514 5290 5594 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05601 7514 5290 5594 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05600 5594 5290 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05599 7514 5296 5231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05598 5232 5231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05597 7514 5231 5232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05596 7514 5231 5232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05595 5232 5231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05594 5583 5586 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05593 5577 5587 5578 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05592 7514 7335 5577 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05591 7514 5584 5587 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05590 5585 5587 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05589 7514 5581 5586 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05588 5579 5582 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05587 7514 5579 5580 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05586 5578 5585 5579 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05585 7335 5578 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05584 7514 5578 7335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05583 5580 5585 5582 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05582 5582 5587 5583 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05581 7514 6266 449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05580 449 4728 484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05579 494 484 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05578 3432 5841 3358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05577 3358 7108 3432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05576 7514 6332 3358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05575 4874 4905 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05574 4872 4906 4899 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05573 7514 5350 4872 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05572 7514 5584 4906 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05571 4904 4906 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05570 7514 5353 4905 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05569 4900 4903 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05568 7514 4900 4873 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05567 4899 4904 4900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05566 5350 4899 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05565 7514 4899 5350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05564 4873 4904 4903 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05563 4903 4906 4874 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05562 7473 7475 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05561 1610 2926 1646 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05560 1646 3135 1611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05559 1611 2949 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05558 1609 2925 1646 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05557 7514 5138 1609 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05556 7514 5882 1610 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05555 1883 1646 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05554 7514 5296 5295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05553 5294 5295 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05552 7514 5295 5294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05551 7514 5295 5294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05550 5294 5295 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05549 7514 5296 5297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05548 5518 5297 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05547 7514 5297 5518 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05546 7514 5297 5518 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05545 5518 5297 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05544 7514 7194 6149 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05543 6148 6149 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05542 7514 6149 6148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05541 7514 6149 6148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05540 6148 6149 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05539 7514 7194 6223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05538 6222 6223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05537 7514 6223 6222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05536 7514 6223 6222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05535 6222 6223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05534 7514 7194 6224 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05533 6622 6224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05532 7514 6224 6622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05531 7514 6224 6622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05530 6622 6224 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05529 7514 7194 6155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05528 6154 6155 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05527 7514 6155 6154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05526 7514 6155 6154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05525 6154 6155 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05524 7514 7194 6230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05523 6229 6230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05522 7514 6230 6229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05521 7514 6230 6229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05520 6229 6230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05519 7514 7194 6232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05518 6231 6232 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05517 7514 6232 6231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05516 7514 6232 6231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05515 6231 6232 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05514 7513 7512 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05513 5860 7335 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05512 4282 4782 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05511 5075 5376 4878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05510 4878 5273 5075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05509 7514 6388 4878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05508 3484 3214 3190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05507 3190 3212 3484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05506 7514 3475 3190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05505 2285 2841 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05504 2286 2836 2285 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05503 7094 7481 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05502 1630 4448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05501 1631 1976 1630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05500 3064 3119 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05499 3667 3266 3064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05498 5345 5992 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05497 5376 5891 5345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05496 6294 7491 6295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05495 6295 7379 6294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05494 7514 7452 6295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05493 6293 6294 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05492 7297 7493 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05491 7514 7493 7331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05490 7514 7494 7296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05489 7329 7330 7297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05488 7296 7331 7329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05487 7315 7329 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05486 7514 7329 7315 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05485 7330 7494 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05484 7514 7194 7125 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05483 7124 7125 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05482 7514 7125 7124 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05481 7514 7125 7124 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05480 7124 7125 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05479 7514 7194 7188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05478 7187 7188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05477 7514 7188 7187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05476 7514 7188 7187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05475 7187 7188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05474 7514 7194 7190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05473 7189 7190 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05472 7514 7190 7189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05471 7514 7190 7189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05470 7189 7190 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05469 7514 7194 7127 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05468 7126 7127 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05467 7514 7127 7126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05466 7514 7127 7126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05465 7126 7127 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05464 7514 7194 7192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05463 7191 7192 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05462 7514 7192 7191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05461 7514 7192 7191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05460 7191 7192 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05459 7514 7194 7195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05458 7193 7195 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05457 7514 7195 7193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05456 7514 7195 7193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05455 7193 7195 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05454 7514 7207 6164 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05453 6163 6164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05452 7514 6164 6163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05451 7514 6164 6163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05450 6163 6164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05449 7499 7510 7502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05448 7498 7509 7499 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05447 7496 7499 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05446 7514 7499 7496 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05445 7506 7507 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05444 7514 7505 7507 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05443 7510 7509 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05442 7514 7508 7509 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05441 7501 7504 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05440 7502 7500 7501 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05439 7504 7509 7506 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05438 7503 7510 7504 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05437 7514 7502 7503 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05436 7514 7496 7497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05435 7497 7500 7498 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05434 7514 6600 6467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05433 7514 6848 6467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05432 6467 6599 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05431 7420 6467 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05430 2963 2970 2964 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05429 2905 2969 2963 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05428 3814 2963 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05427 7514 2963 3814 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05426 2909 2967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05425 7514 2973 2967 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05424 2970 2969 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05423 7514 3263 2969 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05422 2907 2965 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05421 2964 7500 2907 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05420 2965 2969 2909 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05419 2908 2970 2965 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05418 7514 2964 2908 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05417 7514 3814 2906 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05416 2906 7500 2905 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05415 879 2371 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05414 906 1851 879 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05413 340 4376 167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05412 7514 4161 194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05411 167 194 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05410 6220 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05409 6267 6266 6220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05408 7514 7207 6238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05407 6237 6238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05406 7514 6238 6237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05405 7514 6238 6237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05404 6237 6238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05403 7514 7207 6239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05402 6302 6239 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05401 7514 6239 6302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05400 7514 6239 6302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05399 6302 6239 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05398 7514 7207 6171 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05397 6172 6171 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05396 7514 6171 6172 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05395 7514 6171 6172 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05394 6172 6171 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05393 7514 7207 6244 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05392 6243 6244 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05391 7514 6244 6243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05390 7514 6244 6243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05389 6243 6244 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05388 7514 7207 6245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05387 6528 6245 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05386 7514 6245 6528 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05385 7514 6245 6528 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05384 6528 6245 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05383 7514 7207 7134 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05382 7133 7134 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05381 7514 7134 7133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05380 7514 7134 7133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05379 7133 7134 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05378 7514 7207 7198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05377 7197 7198 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05376 7514 7198 7197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05375 7514 7198 7197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05374 7197 7198 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05373 7514 7207 7200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05372 7199 7200 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05371 7514 7200 7199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05370 7514 7200 7199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05369 7199 7200 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05368 7514 6173 4614 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05367 4614 4912 4647 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05366 7514 4912 4648 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05365 4647 4648 4615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05364 4644 4647 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05363 4615 4979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05362 2453 2454 2455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05361 2455 3837 2453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05360 7514 4589 2455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05359 2452 2453 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05358 4439 4448 4438 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05357 4438 4441 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05356 4440 5173 4439 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05355 4594 4446 4440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05354 7221 7491 7181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05353 7181 7379 7221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05352 7514 7489 7181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05351 7219 7221 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05350 6638 7033 6640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05349 6639 6885 6638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05348 6640 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05347 6637 6638 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05346 7514 7032 6639 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05345 6639 7024 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05344 4325 4377 4324 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05343 4324 4447 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05342 4323 4442 4325 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05341 6846 4376 4323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05340 7514 7207 7140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05339 7141 7140 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05338 7514 7140 7141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05337 7514 7140 7141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05336 7141 7140 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05335 7514 7207 7206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05334 7205 7206 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05333 7514 7206 7205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05332 7514 7206 7205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05331 7205 7206 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05330 7514 7207 7209 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05329 7208 7209 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05328 7514 7209 7208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05327 7514 7209 7208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05326 7208 7209 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05325 7514 6739 4753 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05324 5280 4753 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05323 7514 4753 5280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05322 7514 4753 5280 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05321 5280 4753 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05320 2161 2514 2160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05319 2160 2159 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05318 2158 2383 2161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05317 2157 2304 2158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05316 740 819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05315 1022 765 740 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05314 739 1153 1022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05313 7514 905 739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05312 739 1029 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05311 7514 6739 4767 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05310 5296 4767 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05309 7514 4767 5296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05308 7514 4767 5296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05307 5296 4767 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05306 7514 6739 6725 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05305 7194 6725 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05304 7514 6725 7194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05303 7514 6725 7194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05302 7194 6725 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05301 7514 6739 6740 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05300 7207 6740 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05299 7514 6740 7207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05298 7514 6740 7207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05297 7207 6740 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05296 7514 6266 5197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05295 5197 5718 5250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05294 5249 5250 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05293 7514 6473 6216 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05292 6216 6259 6258 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05291 6700 6258 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05290 5026 5066 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05289 5024 5068 5060 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05288 7514 6392 5024 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05287 7514 5594 5068 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05286 5067 5068 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05285 7514 5065 5066 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05284 5061 5064 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05283 7514 5061 5025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05282 5060 5067 5061 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05281 6392 5060 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05280 7514 5060 6392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05279 5025 5067 5064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05278 5064 5068 5026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05277 6631 7491 6630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05276 6630 7379 6631 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05275 7514 7454 6630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05274 4454 4479 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05273 4452 4481 4474 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05272 7514 6025 4452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05271 7514 4638 4481 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05270 4480 4481 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05269 7514 4475 4479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05268 4473 4477 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05267 7514 4473 4453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05266 4474 4480 4473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05265 6025 4474 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05264 7514 4474 6025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05263 4453 4480 4477 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05262 4477 4481 4454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05261 1018 1051 1019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05260 1019 1052 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05259 1017 4448 1018 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05258 6332 1053 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05257 1053 5173 1017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05256 454 893 424 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05255 424 455 454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05254 7514 641 424 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05253 554 454 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05252 6497 6552 6521 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05251 7514 6628 6497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05250 6498 6553 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05249 6521 6551 6498 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05248 7514 6553 6552 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05247 6551 6628 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05246 2932 3957 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05245 7514 2587 2932 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05244 2932 6030 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05243 7514 3958 2932 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05242 6643 6968 6642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05241 6642 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05240 6641 7489 6643 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05239 28 29 470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05238 7514 281 28 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05237 30 325 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05236 470 27 30 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05235 7514 325 29 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05234 27 281 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05233 6504 6968 6503 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05232 6503 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05231 6696 7493 6504 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05230 7514 5234 5194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05229 5194 5233 5236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05228 5235 5236 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05227 2175 4158 2176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05226 2176 2174 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05225 2954 5690 2175 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05224 466 515 465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05223 465 514 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05222 828 1342 466 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05221 7514 2613 2615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05220 2615 2685 2614 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05219 2612 2614 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05218 7514 4732 3685 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05217 3685 3729 3730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05216 4264 3730 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05215 6659 6683 6660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05214 6660 7422 6684 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05213 7514 6882 6659 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05212 6682 6684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05211 6509 6562 6510 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05210 6510 7218 6563 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05209 7514 6641 6509 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05208 6598 6563 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05207 881 1768 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05206 1342 1435 881 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05205 1529 4081 1530 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05204 1530 2033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05203 1528 2103 1529 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05202 1826 7162 1528 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05201 1246 1257 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05200 1858 1258 1246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05199 147 145 461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05198 7514 900 147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05197 148 899 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05196 461 146 148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05195 7514 899 145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05194 146 900 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05193 5456 5454 5455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05192 5455 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05191 5453 5841 5456 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05190 6259 6333 5453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05189 7514 793 531 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05188 721 531 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05187 7514 531 721 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05186 7514 531 721 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05185 721 531 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05184 7514 721 158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05183 4081 158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05182 7514 158 4081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05181 7514 158 4081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05180 4081 158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05179 7514 721 722 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05178 4600 722 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05177 7514 722 4600 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05176 7514 722 4600 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05175 4600 722 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05174 6673 7034 6655 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05173 6654 6731 6673 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05172 6655 7033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05171 6672 6673 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05170 7514 7032 6654 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05169 6654 6817 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05168 7514 3483 3041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05167 3041 3077 3078 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05166 3137 3078 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05165 7514 2811 2770 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05164 2770 2814 2812 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05163 3501 2812 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05162 7356 7512 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05161 7514 7387 7356 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05160 7514 5901 7033 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05159 5901 6047 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05158 7033 6600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05157 4460 4499 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05156 4458 4501 4493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05155 7514 4782 4458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05154 7514 4561 4501 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05153 4500 4501 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05152 7514 4498 4499 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05151 4494 4497 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05150 7514 4494 4459 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05149 4493 4500 4494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05148 4782 4493 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05147 7514 4493 4782 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05146 4459 4500 4497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05145 4497 4501 4460 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05144 151 576 127 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05143 127 470 151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05142 7514 464 127 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05141 126 151 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05140 1535 1572 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05139 2958 2035 1535 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05138 1534 7114 2958 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05137 7514 2174 1534 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05136 1534 1837 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_05135 2330 2687 2329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05134 2329 2684 2331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05133 7514 4000 2330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05132 2328 2331 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05131 2896 3226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05130 3080 3081 2896 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05129 2895 2926 3080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05128 7514 5887 2895 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05127 2894 2925 3080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05126 7514 5274 2894 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05125 6443 7452 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05124 7488 7489 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05123 3992 4215 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05122 4067 4207 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05121 7463 7462 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05120 1014 1976 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05119 1618 1049 1014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05118 2101 2099 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05117 7514 2723 2101 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05116 6090 6576 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05115 6271 6652 6090 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05114 5826 6599 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05113 7514 6406 5826 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05112 5826 5832 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05111 7514 6600 5826 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05110 846 5173 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05109 1112 1908 846 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05108 1113 1112 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05107 1445 1111 1113 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05106 7514 5685 5384 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05105 5384 5467 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05104 5891 5384 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05103 7514 6388 4550 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05102 4550 4912 4552 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05101 7514 4912 4553 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05100 4552 4553 4551 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05099 4635 4552 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05098 4551 5216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05097 2989 3023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05096 2988 6333 2989 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05095 7514 6392 4844 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05094 4844 4912 4913 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05093 7514 4912 4915 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05092 4913 4915 4845 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05091 5065 4913 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05090 4845 5055 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_05089 2843 3484 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05088 2842 3483 2843 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05087 3912 3913 3858 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05086 3858 4360 3912 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05085 7514 6326 3858 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05084 3911 3912 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05083 4322 4600 4321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05082 4321 4603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05081 4320 6266 4322 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05080 4370 7114 4320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05079 5708 5735 5338 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05078 5338 5734 5708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05077 7514 5876 5338 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05076 6384 6393 5883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05075 5883 6394 6384 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05074 7514 5882 5883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05073 7514 4376 757 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05072 757 1449 796 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05071 1384 796 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05070 702 705 3637 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05069 7514 829 702 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05068 704 1034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05067 3637 703 704 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05066 7514 1034 705 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05065 703 829 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05064 4507 6408 4463 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05063 4464 4986 4507 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05062 4463 6407 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05061 4998 4507 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05060 7514 4987 4464 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05059 4464 4984 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05058 4730 6266 4729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05057 4729 4728 4731 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05056 7514 7114 4730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05055 6600 4731 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05054 6989 6990 6939 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05053 6938 7387 6989 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05052 6939 6992 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05051 7343 6989 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05050 7514 6991 6938 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05049 6938 7045 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05048 7514 1304 872 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05047 872 1906 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05046 1575 872 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05045 7514 4784 4815 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05044 4784 4783 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05043 4815 5378 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05042 7514 2256 1949 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05041 1949 2189 1978 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05040 2332 1978 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05039 2458 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05038 4106 2457 2458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05037 7514 2456 4106 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05036 7514 1908 605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05035 605 5173 604 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05034 728 604 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05033 422 450 1023 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05032 7514 1068 422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05031 423 762 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05030 1023 451 423 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05029 7514 762 450 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05028 451 1068 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05027 1407 1575 1408 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05026 1408 1574 1439 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05025 7514 2602 1407 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05024 2040 1439 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_05023 1622 1620 1621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05022 1623 1834 1622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05021 1621 1619 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05020 1974 1622 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05019 7514 5467 1623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05018 1623 1618 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_05017 1800 2037 1801 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05016 1801 1835 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05015 1799 1896 1800 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05014 2333 1836 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_05013 1836 1899 1799 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_05012 2632 2673 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05011 2630 2675 2668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05010 7514 2664 2630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05009 7514 2672 2675 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05008 2674 2675 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_05007 7514 2669 2673 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_05006 2667 2670 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05005 7514 2667 2631 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05004 2668 2674 2667 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05003 2664 2668 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05002 7514 2668 2664 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_05001 2631 2674 2670 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_05000 2670 2675 2632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04999 7514 370 318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04998 318 953 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04997 462 319 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04996 318 372 319 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04995 319 1466 318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04994 700 699 701 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04993 701 698 700 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04992 7514 1341 701 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04991 768 700 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04990 6618 6621 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04989 6588 6619 6616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04988 7514 6617 6588 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04987 7514 6622 6619 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04986 6592 6619 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04985 7514 6620 6621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04984 6589 6590 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04983 7514 6589 6591 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04982 6616 6592 6589 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04981 6617 6616 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04980 7514 6616 6617 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04979 6591 6592 6590 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04978 6590 6619 6618 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04977 5292 5826 5293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04976 5293 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04975 5291 7511 5292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04974 7514 4695 3772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04973 3772 3770 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04972 3769 3773 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04971 3772 4697 3773 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04970 3773 3771 3772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04969 2582 3499 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04968 2583 3135 2582 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04967 2581 2926 2583 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04966 7514 6025 2581 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04965 2580 2925 2583 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04964 7514 5137 2580 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04963 5641 5829 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04962 5676 5675 5641 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04961 1202 1203 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04960 1652 1569 1202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04959 2051 2079 3159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04958 7514 2081 2051 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04957 2052 2082 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04956 3159 2080 2052 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04955 7514 2082 2079 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04954 2080 2081 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04953 7514 6386 6209 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04952 6209 6241 6240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04951 6683 6240 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04950 7514 4411 3627 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04949 3627 3978 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04948 3625 3626 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04947 3627 4413 3626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04946 3626 4838 3627 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04945 5375 5371 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04944 7514 5818 5375 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04943 5375 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04942 7514 5815 5375 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04941 5679 5375 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04940 7514 6957 6212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04939 6212 6247 6248 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04938 6562 6248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04937 7514 4411 3674 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04936 3674 3705 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04935 3701 3703 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04934 3674 4413 3703 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04933 3703 4971 3674 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04932 7514 1661 1976 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04931 1661 2111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04930 1976 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04929 4734 6266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04928 4732 4828 4734 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04927 4733 7162 4732 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04926 7514 4790 4733 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04925 4733 5016 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04924 3166 4987 3165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04923 3165 4984 3166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04922 7514 4986 3165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04921 3326 3166 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04920 7514 6531 6360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04919 6360 6399 6401 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04918 6400 6401 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04917 5683 7334 5633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04916 5633 7383 5683 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04915 7514 7454 5633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04914 7514 4411 3981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04913 3981 4112 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04912 3979 3980 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04911 3981 4413 3980 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04910 3980 5134 3981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04909 7514 6569 6506 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04908 6506 6568 6567 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04907 6532 6567 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04906 6328 7334 6327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04905 6327 7383 6328 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04904 7514 6676 6327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04903 5393 5470 5349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04902 5349 6058 5393 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04901 7514 5693 5349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04900 6346 6374 6372 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04899 7514 6443 6346 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04898 6347 6518 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04897 6372 6371 6347 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04896 7514 6518 6374 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04895 6371 6443 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04894 7514 1577 1005 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04893 1005 2591 1039 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04892 1355 1039 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04891 3990 3992 3991 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04890 3991 4360 3990 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04889 7514 5307 3991 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04888 3989 3990 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04887 7514 987 1385 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04886 987 6266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04885 1385 1168 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04884 7514 3067 3040 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04883 3040 3066 3068 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04882 3074 3068 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04881 7514 1341 1080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04880 1080 1342 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04879 1266 1079 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04878 1080 1270 1079 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04877 1079 1866 1080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04876 2520 2945 2485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04875 2485 2946 2520 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04874 7514 5137 2485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04873 1599 1633 1600 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04872 1600 1636 1635 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04871 7514 1634 1599 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04870 1598 1635 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04869 1604 2008 1603 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04868 1603 1641 1640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04867 7514 1855 1604 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04866 4987 1640 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04865 5488 5751 5489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04864 5489 5537 5538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04863 7514 6955 5488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04862 5539 5538 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04861 7218 7219 7180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04860 7180 7377 7218 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04859 7514 7420 7180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04858 7514 6061 5915 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04857 5915 6652 5916 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04856 7164 5916 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04855 6885 7491 6884 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04854 6884 7379 6885 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04853 7514 7481 6884 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04852 3733 3742 3377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04851 3377 3428 3733 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04850 7514 3427 3377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04849 7514 6337 6339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04848 6339 6338 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04847 7514 7334 6339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04846 4406 4407 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04845 4393 4408 4405 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04844 7514 4642 4393 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04843 7514 4488 4408 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04842 4409 4408 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04841 7514 4765 4407 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04840 4394 4395 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04839 7514 4394 4396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04838 4405 4409 4394 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04837 4642 4405 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04836 7514 4405 4642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04835 4396 4409 4395 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04834 4395 4408 4406 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04833 3739 3993 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04832 3511 3468 3460 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04831 3458 3467 3511 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04830 4148 3511 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04829 7514 3511 4148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04828 3464 3465 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04827 7514 3463 3465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04826 3468 3467 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04825 7514 3466 3467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04824 3459 3462 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04823 3460 7500 3459 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04822 3462 3467 3464 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04821 3461 3468 3462 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04820 7514 3460 3461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04819 7514 4148 3457 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04818 3457 7500 3458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04817 2872 3819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04816 5619 1304 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04815 7287 6991 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04814 2681 2543 2493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04813 2493 2541 2681 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04812 7514 2542 2493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04811 42 162 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04810 41 3120 42 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04809 256 338 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04808 480 2875 256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04807 131 193 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04806 130 2817 131 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04805 6779 6818 6817 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04804 7514 6965 6779 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04803 6780 6869 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04802 6817 6815 6780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04801 7514 6869 6818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04800 6815 6965 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04799 6570 6565 6362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04798 6362 6566 6570 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04797 7514 7453 6362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04796 878 949 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04795 905 951 878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04794 5385 6266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04793 1110 1109 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04792 2541 1111 1110 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04791 134 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04790 295 3346 134 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04789 5628 6968 5627 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04788 5627 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04787 5729 6965 5628 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04786 7514 4934 2471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04785 2471 2813 2472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04784 2688 2472 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04783 6890 7033 6889 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04782 6891 7278 6890 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04781 6889 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04780 6888 6890 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04779 7514 7032 6891 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04778 6891 7274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04777 463 512 430 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04776 429 464 463 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04775 430 571 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04774 566 463 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04773 7514 576 429 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04772 429 470 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04771 948 1809 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04770 949 1271 948 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04769 5988 7334 5900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04768 5900 7383 5988 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04767 7514 7462 5900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04766 6215 6980 6214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04765 6214 6979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04764 6253 7494 6215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04763 1502 1501 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04762 1619 1500 1502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04761 1358 1489 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04760 5734 1694 1358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04759 2725 3160 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04758 3389 3159 2725 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04757 7514 4934 156 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04756 156 6344 188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04755 7514 6344 170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04754 188 170 157 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04753 584 188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04752 157 4979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04751 7514 4161 717 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04750 717 6344 718 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04749 7514 6344 720 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04748 718 720 719 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04747 785 718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04746 719 4834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04745 4249 6166 4250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04744 4250 6165 4249 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04743 7514 5069 4250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04742 399 1168 353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04741 7514 1449 400 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04740 353 400 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04739 4028 4081 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04738 4518 4437 4028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04737 4725 4724 4727 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04736 4727 4726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04735 4819 5178 4725 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04734 7514 1449 436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04733 436 6344 473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04732 7514 6344 474 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04731 473 474 435 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04730 527 473 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04729 435 5274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04728 7514 2111 2046 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04727 2046 6344 2047 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04726 7514 6344 2048 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04725 2047 2048 2045 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04724 2118 2047 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04723 2045 5043 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04722 7278 7491 7279 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04721 7279 7379 7278 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04720 7514 7480 7279 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04719 862 1040 861 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04718 861 1041 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04717 860 4588 862 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04716 1356 4589 860 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04715 1103 1384 1104 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04714 1104 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04713 1102 3820 1103 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04712 1236 2881 1102 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04711 7514 4411 3003 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04710 3003 3001 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04709 3000 3002 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04708 3003 4413 3002 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04707 3002 4852 3003 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04706 7514 3343 2776 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04705 2776 3348 2818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04704 2817 2818 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04703 5764 5801 5763 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04702 5763 6940 5802 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04701 7514 6158 5764 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04700 5952 5802 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04699 7071 7391 7072 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04698 7072 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04697 7070 7113 7071 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04696 7174 7115 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04695 7115 7114 7070 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04694 2482 2926 2512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04693 2512 3135 2483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04692 2483 3500 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04691 2481 2925 2512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04690 7514 5055 2481 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04689 7514 6392 2482 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04688 2510 2512 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04687 458 505 558 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04686 7514 507 458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04685 459 642 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04684 558 506 459 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04683 7514 642 505 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04682 506 507 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04681 7514 1858 1857 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04680 1857 1954 1856 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04679 1855 1856 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04678 1285 1287 1228 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04677 1228 2095 1285 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04676 7514 1284 1228 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04675 1489 1285 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04674 5430 5431 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04673 5424 5433 5425 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04672 7514 5746 5424 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04671 7514 5518 5433 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04670 5432 5433 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04669 7514 5429 5431 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04668 5426 5427 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04667 7514 5426 5428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04666 5425 5432 5426 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04665 5746 5425 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04664 7514 5425 5746 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04663 5428 5432 5427 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04662 5427 5433 5430 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04661 7514 3321 3158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04660 3158 3722 3157 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04659 3156 3157 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04658 7514 2811 2491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04657 2491 2536 2535 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04656 3456 2535 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04655 7514 3502 3196 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04654 3196 3989 3231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04653 3232 3231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04652 2013 2524 2012 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04651 2012 4694 2014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04650 7514 2228 2013 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04649 2139 2014 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04648 1865 2416 1864 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04647 1864 2576 1863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04646 7514 2220 1865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04645 2647 1863 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04644 597 600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04643 592 601 593 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04642 7514 3820 592 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04641 7514 598 601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04640 599 601 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04639 7514 915 600 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04638 595 596 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04637 7514 595 594 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04636 593 599 595 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04635 3820 593 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04634 7514 593 3820 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04633 594 599 596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04632 596 601 597 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04631 2593 4367 2594 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04630 2594 2733 2595 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04629 7514 4724 2593 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04628 2592 2595 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04627 2360 2880 2361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04626 2361 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04625 2359 4446 2360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04624 2536 2393 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04623 2393 2881 2359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04622 247 268 1144 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04621 7514 266 247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04620 248 1680 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04619 1144 265 248 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04618 7514 1680 268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04617 265 266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04616 2996 3481 2997 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04615 2997 4695 2996 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04614 7514 3077 2997 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04613 3079 2996 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04612 1128 3814 1129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04611 1129 2174 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04610 1127 4158 1128 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04609 1732 1158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04608 1158 5690 1127 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04607 2324 2543 2323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04606 2323 2541 2324 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04605 7514 2322 2323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04604 3023 2324 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04603 139 173 1465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04602 7514 1332 139 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04601 140 312 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04600 1465 174 140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04599 7514 312 173 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04598 174 1332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04597 3252 4569 3200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04596 3200 3655 3252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04595 7514 3659 3200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04594 3348 3252 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04593 4609 4637 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04592 4607 4640 4630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04591 7514 6388 4607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04590 7514 4638 4640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04589 4639 4640 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04588 7514 4635 4637 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04587 4632 4633 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04586 7514 4632 4608 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04585 4630 4639 4632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04584 6388 4630 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04583 7514 4630 6388 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04582 4608 4639 4633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04581 4633 4640 4609 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04580 4923 5376 4880 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04579 4880 5273 4923 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04578 7514 6173 4880 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04577 6761 6169 6070 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04576 6070 6168 6761 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04575 7514 6125 6070 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04574 7514 5377 5381 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04573 5381 6910 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04572 7514 5378 5381 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04571 7514 6991 6915 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04570 7514 7387 6915 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04569 6915 7512 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04568 6914 6915 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04567 7514 4852 3018 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04566 3018 3667 3111 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04565 7514 3667 3113 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04564 3111 3113 3019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04563 3108 3111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04562 3019 3109 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_04561 2457 5467 2206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04560 2206 2256 2457 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04559 7514 2257 2206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04558 7469 7472 7470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04557 7514 7473 7469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04556 7468 7471 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04555 7470 7467 7468 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04554 7514 7471 7472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04553 7467 7473 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04552 5898 6980 5899 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04551 5899 6979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04550 5897 7493 5898 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04549 5315 7108 5316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04548 5314 5840 5315 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04547 5316 5842 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04546 5876 5315 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04545 7514 5841 5314 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04544 5314 6133 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04543 7101 7280 7064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04542 7064 7428 7101 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04541 7514 7493 7064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04540 7514 76 181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04539 76 3546 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04538 181 2134 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04537 1796 2813 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04536 1893 2536 1796 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04535 6055 6266 6054 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04534 6054 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04533 6194 7114 6055 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04532 4853 4852 4854 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04531 4854 5369 4853 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04530 7514 5226 4854 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04529 5967 4853 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04528 7514 4674 4624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04527 4624 4673 4675 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04526 6405 4675 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04525 4564 4566 4567 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04524 4565 4986 4564 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04523 4567 5085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04522 4809 4564 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04521 7514 4987 4565 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04520 4565 4984 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04519 3502 3501 3503 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04518 3503 4669 3502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04517 7514 3500 3503 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04516 3322 3501 3323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04515 3323 4669 3322 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04514 7514 3645 3323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04513 7514 6056 5634 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04512 5634 6773 5694 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04511 5693 5694 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04510 1613 1700 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04509 1750 1968 1613 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04508 1612 1967 1750 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04507 7514 5735 1612 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04506 1612 5734 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04505 2841 3214 2840 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04504 2840 3212 2841 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04503 7514 6617 2840 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04502 7514 3352 3114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04501 3114 4158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04500 3428 3114 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04499 1948 2880 1947 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04498 1947 2591 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04497 1946 4446 1948 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04496 2257 2881 1946 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04495 7514 1732 1735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04494 1735 1954 1734 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04493 1733 1734 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04492 7514 3266 3038 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04491 3038 3119 3039 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04490 3037 3039 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04489 2476 2504 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04488 3407 2505 2476 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04487 2475 3138 3407 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04486 7514 2502 2475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04485 2474 2789 3407 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04484 7514 2794 2474 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04483 7514 2379 2507 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04482 2379 2520 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04481 2507 2986 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04480 7514 6570 6507 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04479 6507 6572 6571 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04478 6644 6571 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04477 7514 4732 4621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04476 4621 5093 4668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04475 4667 4668 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04474 6937 6980 6936 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04473 6936 6979 6978 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04472 7514 7475 6937 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04471 6954 6978 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04470 6669 6707 6668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04469 6668 7234 6709 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04468 7514 6708 6669 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04467 6902 6709 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04466 7514 7283 7284 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04465 7427 7284 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04464 7514 7284 7427 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04463 7514 7284 7427 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04462 7427 7284 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04461 7514 7427 7429 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04460 7428 7429 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04459 7514 7429 7428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04458 7514 7429 7428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04457 7428 7429 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04456 7514 7427 7380 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04455 7379 7380 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04454 7514 7380 7379 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04453 7514 7380 7379 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04452 7379 7380 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04451 1766 1764 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04450 3178 1765 1766 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04449 1763 7114 3178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04448 7514 2174 1763 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04447 1763 1837 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04446 772 3081 742 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04445 742 1187 772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04444 7514 771 742 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04443 824 772 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04442 1208 1365 1207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04441 1207 1501 1208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04440 7514 1500 1207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04439 2179 1208 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04438 1918 1955 6166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04437 7514 1952 1918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04436 1919 1954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04435 6166 1951 1919 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04434 7514 1954 1955 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04433 1951 1952 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04432 4017 4062 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04431 4015 4064 4057 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04430 7514 4069 4015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04429 7514 4561 4064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04428 4063 4064 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04427 7514 4059 4062 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04426 4058 4060 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04425 7514 4058 4016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04424 4057 4063 4058 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04423 4069 4057 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04422 7514 4057 4069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04421 4016 4063 4060 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04420 4060 4064 4017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04419 7514 6393 6967 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04418 6967 6315 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04417 7514 6394 6967 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04416 4988 4985 4990 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04415 4989 4986 4988 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04414 4990 5085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04413 5879 4988 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04412 7514 4987 4989 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04411 4989 4984 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04410 3505 3506 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04409 3452 3508 3504 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04408 7514 3727 3452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04407 7514 3581 3508 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04406 3507 3508 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04405 7514 3648 3506 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04404 3453 3455 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04403 7514 3453 3454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04402 3504 3507 3453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04401 3727 3504 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04400 7514 3504 3727 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04399 3454 3507 3455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04398 3455 3508 3505 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04397 7098 7144 7062 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04396 7062 7372 7098 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04395 7514 7420 7062 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04394 2881 2111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04393 4000 2686 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04392 3742 3820 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04391 1090 3023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04390 1271 3814 1090 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04389 5917 6061 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04388 5467 7162 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04387 6019 6968 6018 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04386 6018 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04385 6017 7335 6019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04384 2744 6133 2745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04383 2745 5994 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04382 2743 4934 2744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04381 6122 7034 6080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04380 6079 6380 6122 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04379 6080 7033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04378 6096 6122 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04377 7514 7032 6079 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04376 6079 6521 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04375 6476 6474 6475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04374 6475 6894 6476 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04373 7514 6901 6475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04372 7514 4724 4465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04371 4465 4726 4509 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04370 4582 4509 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04369 471 3081 433 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04368 433 1085 471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04367 7514 831 433 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04366 654 471 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04365 1375 4158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04364 1373 3427 1375 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04363 1374 1371 1373 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04362 7514 5467 1374 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04361 1374 1372 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04360 627 4081 626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04359 626 1292 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04358 625 963 627 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04357 1040 5841 625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04356 7514 3135 1642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04355 7514 1736 1642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04354 1642 1959 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04353 1684 1642 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04352 2914 3636 2913 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04351 2913 2932 2933 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04350 7514 3637 2914 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04349 2999 2933 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04348 380 3081 350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04347 350 1085 380 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04346 7514 775 350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04345 469 380 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04344 7311 7491 7293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04343 7293 7379 7311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04342 7514 7475 7293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04341 7514 2085 2053 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04340 2053 2140 2084 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04339 2217 2084 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04338 7514 2738 2740 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04337 2740 2739 2742 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04336 2741 2742 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04335 2338 2602 2132 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04334 7514 4161 2194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04333 2132 2194 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04332 5470 7388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04331 3500 4861 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04330 3644 4716 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04329 693 1145 692 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04328 692 1029 694 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04327 7514 829 693 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04326 691 694 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04325 7514 6701 6703 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04324 6701 6700 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04323 6703 6841 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04322 2078 6980 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04321 2319 6979 2078 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04320 2077 2322 2319 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04319 7514 2543 2077 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04318 2077 2541 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04317 3499 4502 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04316 2949 4504 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04315 6778 6812 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04314 6776 6814 6806 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04313 7514 6804 6776 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04312 7514 7189 6814 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04311 6813 6814 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04310 7514 6811 6812 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04309 6807 6810 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04308 7514 6807 6777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04307 6806 6813 6807 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04306 6804 6806 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04305 7514 6806 6804 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04304 6777 6813 6810 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04303 6810 6814 6778 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04302 6123 7034 6082 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04301 6081 6124 6123 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04300 6082 7033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04299 6099 6123 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04298 7514 7032 6081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04297 6081 6678 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_04296 283 653 255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04295 255 654 283 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04294 7514 777 255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04293 5648 5841 5649 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04292 5649 5691 5692 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04291 7514 5690 5648 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04290 6337 5692 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04289 2893 3644 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04288 2922 3135 2893 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04287 2892 2926 2922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04286 7514 6388 2892 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04285 2891 2925 2922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04284 7514 5216 2891 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04283 2885 6342 2886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04282 2886 2951 2885 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04281 7514 2884 2886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04280 2887 2885 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04279 4404 5826 4403 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04278 4403 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04277 4755 4959 4404 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04276 5896 6107 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04275 5895 6180 5896 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04274 5436 5435 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04273 7514 5818 5436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04272 5436 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04271 7514 5815 5436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04270 5434 5436 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04269 1666 3081 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04268 1727 3646 1666 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04267 4843 4841 4842 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04266 4842 5369 4843 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04265 7514 5226 4842 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04264 5413 4843 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04263 5234 5376 5030 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04262 5030 5273 5234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04261 7514 5882 5030 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04260 1476 1686 1475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04259 1475 1473 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04258 1474 1550 1476 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04257 3024 3170 3025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04256 3025 3917 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04255 3347 5225 3024 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04254 519 653 490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04253 490 654 519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04252 7514 833 490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04251 706 519 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04250 4327 4368 4328 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04249 4328 5085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04248 4326 4367 4327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04247 4401 4357 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_04246 4357 4985 4326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04245 7514 2541 1410 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04244 1410 2543 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04243 1444 1448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04242 1410 2179 1448 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04241 1448 1445 1410 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04240 234 237 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04239 229 238 230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04238 7514 1304 229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04237 7514 669 238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04236 236 238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04235 7514 233 237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04234 231 235 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04233 7514 231 232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04232 230 236 231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04231 1304 230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04230 7514 230 1304 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04229 232 236 235 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04228 235 238 234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04227 2429 2661 2297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04226 2297 2658 2429 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04225 7514 2502 2297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04224 2421 2507 2423 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04223 2423 3769 2422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04222 7514 2508 2421 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04221 3549 2422 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04220 2771 2813 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04219 2869 2814 2771 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04218 7514 2872 2869 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04217 7514 6253 5933 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04216 5933 5984 5983 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04215 5982 5983 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04214 7514 6846 5347 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04213 5347 5385 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04212 5386 5389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04211 5347 5387 5389 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04210 5389 6845 5347 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_04209 5645 5683 5644 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04208 5644 5681 5682 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04207 7514 6185 5645 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04206 5810 5682 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04205 5614 5617 5615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04204 5615 5616 5614 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04203 7514 5889 5615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04202 6893 5614 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04201 3483 3418 2897 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04200 2897 2929 3483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04199 7514 5887 2897 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04198 6015 6014 6016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04197 6016 6375 6015 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04196 7514 7420 6016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04195 1536 1575 1537 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04194 1537 1574 1576 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04193 7514 2255 1536 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04192 2042 1576 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04191 3540 3734 3598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04190 3598 3733 3541 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04189 3541 3732 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04188 3539 3920 3598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04187 7514 4077 3539 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04186 7514 3967 3540 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04185 6980 3598 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04184 143 176 1332 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04183 7514 1413 143 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04182 144 1736 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04181 1332 177 144 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04180 7514 1736 176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04179 177 1413 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04178 4856 4858 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04177 4811 4860 4855 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04176 7514 5160 4811 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04175 7514 5531 4860 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04174 4859 4860 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04173 7514 4857 4858 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04172 4812 4813 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04171 7514 4812 4814 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04170 4855 4859 4812 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04169 5160 4855 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04168 7514 4855 5160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04167 4814 4859 4813 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04166 4813 4860 4856 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04165 5181 5188 5182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04164 5180 5189 5181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04163 7390 5181 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04162 7514 5181 7390 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04161 5186 5187 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04160 7514 5331 5187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04159 5188 5189 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04158 7514 5554 5189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04157 5183 5185 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04156 5182 7500 5183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04155 5185 5189 5186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04154 5184 5188 5185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04153 7514 5182 5184 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04152 7514 7390 5179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04151 5179 7500 5180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04150 5751 7334 5750 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04149 5750 7383 5751 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04148 7514 6628 5750 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04147 7514 6134 6114 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04146 6134 6533 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04145 6114 6538 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04144 7514 2340 2813 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04143 2340 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04142 2813 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04141 1859 1954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04140 2009 1858 1859 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04139 7514 2093 4986 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04138 4986 2090 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04137 7514 2091 4986 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04136 21 22 900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04135 7514 272 21 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04134 20 181 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04133 900 19 20 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04132 7514 181 22 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04131 19 272 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04130 6513 7286 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04129 6533 7384 6513 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04128 2866 2953 2867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04127 2867 2865 2866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04126 7514 3108 2867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04125 1525 1567 1526 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04124 1526 3160 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04123 1749 3159 1525 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04122 2919 2954 2918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04121 2918 3179 2955 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04120 7514 2995 2919 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04119 2953 2955 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04118 5719 5718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04117 6907 6133 5719 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04116 3509 4600 3510 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04115 3510 4603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04114 4367 7108 3509 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04113 4999 5834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04112 5256 4998 4999 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04111 5630 6968 5629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04110 5629 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04109 5807 6628 5630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04108 6312 6310 6311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04107 6311 7212 6313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04106 7514 6831 6312 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04105 6309 6313 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04104 6635 6633 6634 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04103 6634 6948 6636 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04102 7514 6741 6635 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04101 6632 6636 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04100 7514 4923 4739 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04099 4739 4771 4772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04098 5079 4772 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04097 1209 1236 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04096 1235 1441 1209 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04095 7514 1440 1235 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04094 6407 1235 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04093 7430 7227 7182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04092 7182 7228 7430 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04091 7514 7489 7182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04090 7514 6194 6197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04089 6197 6195 6196 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04088 6193 6196 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04087 5932 6037 5931 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04086 5931 6322 5980 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04085 7514 6391 5932 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04084 6032 5980 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04083 5206 5252 5205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04082 5205 5757 5253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04081 7514 5386 5206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04080 5251 5253 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_04079 999 1700 998 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04078 998 1968 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04077 997 1435 999 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04076 1851 1688 997 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04075 1701 2103 1650 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04074 1650 4726 1701 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04073 7514 4773 1650 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04072 1700 1701 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04071 1512 4446 1513 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04070 1513 1775 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04069 1511 1915 1512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04068 4597 3742 1511 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04067 323 571 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04066 823 512 323 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04065 322 464 823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04064 7514 576 322 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04063 322 470 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_04062 568 3081 569 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04061 569 1187 568 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04060 7514 771 569 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04059 5163 5160 5162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04058 5162 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04057 5161 5841 5163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04056 5608 6333 5161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04055 7514 7168 6911 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04054 6911 6912 6913 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04053 6910 6913 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04052 7514 6412 6990 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04051 6412 6410 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04050 6990 6652 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04049 7514 3563 3488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04048 3488 3562 3489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04047 3487 3489 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04046 3238 3501 2902 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04045 2902 4669 3238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04044 7514 3646 2902 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04043 7514 2133 1923 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04042 1923 2424 1960 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04041 1959 1960 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04040 5930 5977 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04039 5928 5978 5971 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04038 7514 5969 5928 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04037 7514 6693 5978 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04036 5979 5978 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_04035 7514 5974 5977 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_04034 5972 5976 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04033 7514 5972 5929 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04032 5971 5979 5972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04031 5969 5971 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04030 7514 5971 5969 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04029 5929 5979 5976 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04028 5976 5978 5930 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04027 7514 2861 2863 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04026 2863 3233 2864 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04025 2862 2864 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04024 7514 1049 871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04023 871 1976 916 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04022 1628 916 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04021 555 559 3632 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04020 7514 554 555 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04019 557 558 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04018 3632 556 557 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04017 7514 558 559 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04016 556 554 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_04015 1634 1728 612 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04014 612 937 1634 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04013 7514 1681 612 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04012 7514 1258 1181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04011 1181 1257 1220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04010 1952 1220 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04009 7263 7261 7262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04008 7262 7411 7263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04007 7514 7420 7262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04006 6886 7280 6887 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04005 6887 7428 6886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04004 7514 7466 6887 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_04003 4144 4143 4145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04002 4145 4360 4144 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04001 7514 6646 4145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_04000 4142 4144 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03999 4186 5001 4187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03998 4187 5718 4229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03997 7514 4934 4186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03996 4228 4229 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03995 7514 4446 1777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03994 1777 1775 1776 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03993 1911 1776 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03992 54 90 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03991 52 92 84 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03990 7514 286 52 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03989 7514 598 92 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03988 91 92 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03987 7514 656 90 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03986 86 87 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03985 7514 86 53 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03984 84 91 86 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03983 286 84 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03982 7514 84 286 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03981 53 91 87 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03980 87 92 54 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03979 4866 5171 4868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03978 4868 5172 4867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03977 7514 5173 4866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03976 5840 4867 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03975 4871 5470 4870 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03974 4870 5695 4871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03973 7514 6344 4870 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03972 4869 4871 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03971 2956 2537 2358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03970 2358 2390 2956 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03969 7514 7162 2358 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03968 43 65 1681 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03967 7514 262 43 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03966 44 1852 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03965 1681 63 44 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03964 7514 1852 65 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03963 63 262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03962 3354 3352 3353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03961 3353 4673 3354 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03960 7514 4148 3353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03959 3351 3354 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03958 1305 1579 1243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03957 1243 1765 1305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03956 7514 1304 1243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03955 1508 1305 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03954 4363 4361 4318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03953 4318 4360 4363 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03952 7514 6469 4318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03951 4359 4363 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03950 3538 6979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03949 4589 6980 3538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03948 5458 5457 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03947 5617 6333 5458 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03946 1029 696 697 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03945 697 767 1029 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03944 7514 695 697 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03943 3144 3142 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03942 3563 3143 3144 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03941 747 778 746 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03940 746 777 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03939 909 776 747 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03938 3523 3633 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03937 3870 3632 3523 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03936 6076 6133 6075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03935 6075 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03934 6112 7114 6076 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03933 6988 6342 6198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03932 6198 6340 6988 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03931 7514 6713 6198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03930 5192 5826 5191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03929 5191 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03928 5286 7495 5192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03927 5151 6451 5150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03926 5150 5235 5152 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03925 7514 5434 5151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03924 5230 5152 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03923 1755 2315 1754 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03922 1754 1825 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03921 2502 1826 1755 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03920 1663 1684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03919 1682 1813 1663 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03918 1662 1679 1682 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03917 7514 1680 1662 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03916 1662 1681 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03915 6364 6843 6365 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03914 6365 6405 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03913 6363 6768 6364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03912 6406 6907 6363 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03911 1921 2926 1957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03910 1957 3135 1922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03909 1922 3646 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03908 1920 2925 1957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03907 7514 4834 1920 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03906 7514 6175 1921 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03905 2222 1957 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03904 5781 6407 5782 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03903 5782 5837 5838 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03902 7514 6408 5781 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03901 6048 5838 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03900 1086 2435 1087 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03899 1087 2853 1086 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03898 7514 2133 1087 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03897 1085 1086 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03896 817 3625 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03895 1334 2290 817 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03894 816 3546 1334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03893 7514 3549 816 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03892 816 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03891 2682 5467 2640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03890 2640 2681 2682 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03889 7514 2743 2640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03888 3029 2682 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03887 3902 3910 3903 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03886 3853 3909 3902 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03885 4718 3902 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03884 7514 3902 4718 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03883 3857 3908 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03882 7514 3905 3908 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03881 3910 3909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03880 7514 4277 3909 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03879 3855 3907 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03878 3903 5100 3855 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03877 3907 3909 3857 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03876 3856 3910 3907 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03875 7514 3903 3856 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03874 7514 4718 3854 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03873 3854 5100 3853 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03872 3743 3744 3693 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03871 3693 5000 3743 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03870 7514 4378 3693 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03869 7145 7280 7146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03868 7146 7428 7145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03867 7514 7480 7146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03866 7144 7145 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03865 2351 2926 2377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03864 2377 3135 2350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03863 2350 3645 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03862 2349 2925 2377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03861 7514 5043 2349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03860 7514 6035 2351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03859 2433 2377 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03858 7514 2536 2066 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03857 2066 2813 2110 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03856 2109 2110 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03855 7514 5001 610 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03854 610 4728 611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03853 609 611 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03852 4625 5385 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03851 4676 5619 4625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03850 7514 6846 4676 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03849 1792 2101 1791 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03848 1791 2241 1824 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03847 7514 2165 1792 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03846 1823 1824 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03845 7392 7409 7411 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03844 7514 7463 7392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03843 7393 7413 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03842 7411 7410 7393 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03841 7514 7413 7409 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03840 7410 7463 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03839 4129 4130 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03838 4125 4131 4124 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03837 7514 4207 4125 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03836 7514 4561 4131 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03835 4132 4131 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03834 7514 4206 4130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03833 4126 4128 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03832 7514 4126 4127 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03831 4124 4132 4126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03830 4207 4124 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03829 7514 4124 4207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03828 4127 4132 4128 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03827 4128 4131 4129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03826 1743 3004 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03825 1741 1740 1743 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03824 1742 3546 1741 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03823 7514 1823 1742 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03822 1742 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03821 1432 2023 1401 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03820 1401 1823 1432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03819 7514 1431 1401 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03818 1747 1432 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03817 4065 4067 4021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03816 4021 4360 4065 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03815 7514 5982 4021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03814 4066 4065 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03813 5877 6030 5878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03812 5878 6029 5877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03811 7514 5876 5878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03810 2643 2687 2644 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03809 2644 2688 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03808 2972 2686 2643 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03807 7514 5499 5502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03806 5499 5498 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03805 5502 5500 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03804 7271 7272 7270 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03803 7514 7424 7271 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03802 7269 7474 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03801 7270 7268 7269 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03800 7514 7474 7272 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03799 7268 7424 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03798 4524 4676 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03797 7514 4604 4524 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03796 4524 4790 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03795 7514 4679 4524 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03794 4918 4916 4877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03793 4877 5369 4918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03792 7514 5226 4877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03791 5662 4918 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03790 7337 7341 7338 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03789 7303 7342 7337 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03788 7387 7337 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03787 7514 7337 7387 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03786 7306 7340 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03785 7514 7343 7340 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03784 7341 7342 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03783 7514 7508 7342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03782 7304 7339 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03781 7338 7500 7304 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03780 7339 7342 7306 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03779 7305 7341 7339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03778 7514 7338 7305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03777 7514 7387 7302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03776 7302 7500 7303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03775 128 2016 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03774 281 3546 128 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03773 6181 6565 6182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03772 6182 6566 6181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03771 7514 7462 6182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03770 2706 2705 2709 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03769 2709 2708 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03768 2707 2795 2706 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03767 6068 6968 6069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03766 6069 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03765 6102 6676 6068 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03764 619 1732 618 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03763 618 1029 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03762 642 951 619 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03761 7514 731 730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03760 7514 729 730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03759 730 728 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03758 790 730 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03757 687 942 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03756 1680 939 687 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03755 686 685 1680 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03754 7514 1021 686 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03753 686 1022 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03752 4884 5043 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03751 5083 5832 4884 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03750 7514 4929 5083 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03749 4153 4600 4155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03748 4155 4603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03747 4154 6266 4153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03746 5832 4152 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03745 4152 7114 4154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03744 155 653 129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03743 129 654 155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03742 7514 777 129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03741 468 155 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03740 1523 1883 1524 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03739 1524 1565 1566 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03738 7514 1699 1523 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03737 1695 1566 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03736 7130 7132 7129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03735 7514 7454 7130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03734 7131 7460 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03733 7129 7128 7131 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03732 7514 7460 7132 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03731 7128 7454 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03730 7514 5841 5017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03729 5017 5691 5018 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03728 5016 5018 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03727 2326 5467 2327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03726 2327 2454 2326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03725 7514 2325 2327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03724 2730 2326 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03723 1697 1823 1668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03722 1667 2164 1697 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03721 1668 2023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03720 1694 1697 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03719 7514 1695 1667 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03718 1667 1819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03717 123 142 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03716 119 125 141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03715 7514 3868 119 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03714 7514 368 125 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03713 124 125 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03712 7514 3876 142 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03711 120 121 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03710 7514 120 122 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03709 141 124 120 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03708 3868 141 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03707 7514 141 3868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03706 122 124 121 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03705 121 125 123 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03704 2633 2676 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03703 2945 2956 2633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03702 5635 5659 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03701 6119 5655 5635 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03700 4580 4726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03699 4579 4724 4580 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03698 7514 3727 3647 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03697 3647 4577 3650 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03696 7514 4577 3652 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03695 3650 3652 3651 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03694 3648 3650 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03693 3651 3649 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03692 7514 4782 4315 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03691 4315 4577 4356 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03690 7514 4577 4337 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03689 4356 4337 4316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03688 4498 4356 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03687 4316 5127 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03686 7514 4069 3802 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03685 3802 4577 3803 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03684 7514 4577 3805 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03683 3803 3805 3801 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03682 4059 3803 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03681 3801 3804 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03680 3968 4079 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03679 3967 3966 3968 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03678 4470 6846 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03677 7514 4593 4470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03676 4470 4594 5377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03675 5377 5385 4470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03674 5709 5805 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03673 5870 5708 5709 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03672 7514 4207 4179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03671 4179 4577 4210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03670 7514 4577 4212 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03669 4210 4212 4180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03668 4206 4210 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03667 4180 4211 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03666 3189 4934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03665 3837 4158 3189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03664 7514 4695 4700 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03663 4700 4696 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03662 4694 4699 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03661 4700 4697 4699 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03660 4699 4698 4700 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_03659 7514 2596 2598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03658 2598 5128 2600 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03657 7514 5128 2601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03656 2600 2601 2599 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03655 2597 2600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03654 2599 3389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03653 3198 4070 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03652 3239 3238 3198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03651 6370 7391 6369 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03650 6369 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03649 6576 7162 6370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03648 7505 7113 7069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03647 7069 7163 7505 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03646 7514 7111 7069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03645 7019 7033 7021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03644 7020 7311 7019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03643 7021 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03642 7018 7019 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03641 7514 7032 7020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03640 7020 7366 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03639 351 3352 352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03638 352 3820 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03637 481 4376 351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03636 460 462 428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03635 427 511 460 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03634 428 1032 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03633 695 460 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03632 7514 1466 427 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03631 427 461 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03630 4444 4447 4443 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03629 4443 4448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03628 4445 4442 4444 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03627 5387 4934 4445 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03626 1025 1021 991 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03625 991 1022 1025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03624 7514 1023 991 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03623 3982 3955 3949 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03622 3947 3956 3982 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03621 4431 3982 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03620 7514 3982 4431 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03619 3952 3954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03618 7514 3953 3954 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03617 3955 3956 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03616 7514 4488 3956 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03615 3948 3951 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03614 3949 7500 3948 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03613 3951 3956 3952 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03612 3950 3955 3951 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03611 7514 3949 3950 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03610 7514 4431 3946 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03609 3946 7500 3947 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03608 6464 5884 5886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03607 5886 5885 6464 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03606 7514 6315 5886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03605 4079 4934 4027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03604 7514 4158 4080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03603 4027 4080 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03602 7514 5000 1360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03601 1360 1577 1359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03600 2789 1359 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03599 57 99 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03598 55 101 93 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03597 7514 190 55 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03596 7514 669 101 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03595 100 101 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03594 7514 130 99 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03593 95 96 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03592 7514 95 56 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03591 93 100 95 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03590 190 93 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03589 7514 93 190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03588 56 100 96 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03587 96 101 57 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03586 7514 3009 3011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03585 3011 3720 3010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03584 3077 3010 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03583 7514 1569 1403 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03582 1403 1568 1434 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03581 3212 1434 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03580 1545 1727 1515 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03579 1514 3546 1545 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03578 1515 3979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03577 1543 1545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03576 7514 2139 1514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03575 1514 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03574 7514 6042 5610 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03573 5610 5608 5609 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03572 6039 5609 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03571 5153 4991 4992 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03570 4992 5381 5153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03569 7514 6957 4992 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03568 3334 3342 3335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03567 3331 3341 3334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03566 4156 3334 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03565 7514 3334 4156 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03564 3339 3340 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03563 7514 3338 3340 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03562 3342 3341 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03561 7514 3466 3341 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03560 3333 3337 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03559 3335 5100 3333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03558 3337 3341 3339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03557 3336 3342 3337 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03556 7514 3335 3336 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03555 7514 4156 3332 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03554 3332 5100 3331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03553 6948 6969 6922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03552 6922 7092 6948 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03551 7514 7420 6922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03550 882 910 883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03549 883 1341 911 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03548 7514 909 882 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03547 3958 911 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03546 7514 7384 7158 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03545 7158 7353 7159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03544 7228 7159 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03543 3463 3655 3061 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03542 3061 3116 3463 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03541 7514 3183 3061 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03540 4723 4834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03539 4927 5832 4723 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03538 7514 4722 4927 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03537 2231 2661 2200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03536 2200 2658 2231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03535 7514 2510 2200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03534 2229 2231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03533 1503 2543 1504 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03532 1504 2541 1503 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03531 7514 1628 1504 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03530 2174 1503 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03529 3998 3997 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03528 5537 4228 3998 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03527 3996 4156 5537 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03526 7514 4149 3996 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03525 3996 5909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03524 2462 2880 2461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03523 2461 2591 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03522 2460 4446 2462 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03521 2814 2459 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03520 2459 2881 2460 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03519 1705 2543 1655 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03518 1655 2541 1705 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03517 7514 2035 1655 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03516 1880 1705 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03515 7483 7487 7484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03514 7514 7489 7483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03513 7485 7486 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03512 7484 7482 7485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03511 7514 7486 7487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03510 7482 7489 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03509 1480 3023 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03508 2164 2392 1480 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03507 7320 7334 7300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03506 7300 7383 7320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03505 7514 7335 7300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03504 1186 1422 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03503 1337 1474 1186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03502 7514 2647 3411 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03501 3411 2648 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03500 7514 2655 3411 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03499 6378 6625 6349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03498 6349 6942 6378 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03497 7514 7420 6349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03496 3827 3834 3828 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03495 3824 3835 3827 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03494 3993 3827 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03493 7514 3827 3993 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03492 3832 3833 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03491 7514 3830 3833 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03490 3834 3835 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03489 7514 4305 3835 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03488 3826 3831 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03487 3828 7500 3826 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03486 3831 3835 3832 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03485 3829 3834 3831 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03484 7514 3828 3829 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03483 7514 3993 3825 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03482 3825 7500 3824 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03481 6651 6610 6603 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03480 6602 6612 6651 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03479 6652 6651 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03478 7514 6651 6652 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03477 6607 6609 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03476 7514 6608 6609 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03475 6610 6612 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03474 7514 6611 6612 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03473 6604 6606 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03472 6603 7500 6604 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03471 6606 6612 6607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03470 6605 6610 6606 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03469 7514 6603 6605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03468 7514 6652 6601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03467 6601 7500 6602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03466 3180 3178 3182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03465 3182 3181 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03464 3184 3179 3180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03463 6241 6393 6026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03462 6026 6394 6241 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03461 7514 6025 6026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03460 849 1114 848 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03459 848 1632 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03458 847 875 849 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03457 425 1145 426 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03456 426 1029 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03455 893 829 425 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03454 1426 1682 1396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03453 1396 1479 1426 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03452 7514 1556 1396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03451 2465 2398 2365 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03450 2365 2813 2465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03449 7514 2536 2365 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03448 5745 6600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03447 7514 6599 5745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03446 5745 6406 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03445 7514 5832 5745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03444 5818 5745 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03443 2772 3023 2773 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03442 2773 2816 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03441 3179 7114 2772 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03440 5140 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03439 5418 7286 5140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03438 5139 5138 5418 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03437 7514 5275 5139 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03436 5139 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03435 1939 2033 1938 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03434 1938 1970 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03433 1937 4600 1939 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03432 2171 6333 1937 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03431 6038 6407 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03430 6125 6408 6038 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03429 4744 4782 4743 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03428 4743 5718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03427 4742 5001 4744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03426 6707 4934 4742 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03425 5937 6704 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03424 5991 6027 5937 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03423 4779 6894 4741 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03422 4741 4777 4779 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03421 7514 5242 4741 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03420 2586 3500 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03419 2708 3135 2586 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03418 2585 2926 2708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03417 7514 6392 2585 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03416 2584 2925 2708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03415 7514 5055 2584 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03414 7514 7389 7391 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03413 7389 7388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03412 7391 7390 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03411 7514 3742 1916 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03410 1916 1915 1917 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03409 1914 1917 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03408 851 891 6316 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03407 7514 893 851 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03406 853 894 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03405 6316 892 853 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03404 7514 894 891 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03403 892 893 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03402 7514 7494 7401 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03401 7401 7493 7426 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03400 7486 7426 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03399 6511 7286 6512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03398 6512 7164 6564 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03397 7514 7113 6511 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03396 6529 6564 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03395 5178 7388 5177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03394 5177 7390 5178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03393 7514 7384 5177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03392 4746 5620 4745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03391 4745 5387 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03390 4828 4789 4746 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03389 2500 3129 2473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03388 2473 4695 2500 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03387 7514 2841 2473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03386 2785 2500 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03385 7514 7287 7050 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03384 7050 7236 7051 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03383 7049 7051 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03382 2064 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03381 7514 2814 2063 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03380 2104 2536 2064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03379 2063 2103 2104 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03378 7514 2504 2344 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03377 2344 2418 2370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03376 3071 2370 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03375 5483 5529 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03374 5481 5533 5524 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03373 7514 5523 5481 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03372 7514 5531 5533 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03371 5532 5533 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03370 7514 5676 5529 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03369 5526 5528 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03368 7514 5526 5482 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03367 5524 5532 5526 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03366 5523 5524 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03365 7514 5524 5523 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03364 5482 5532 5528 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03363 5528 5533 5483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03362 7514 7108 6767 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03361 6767 7109 6766 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03360 7227 6766 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03359 5337 5360 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03358 5335 5362 5355 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03357 7514 7495 5335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03356 7514 5594 5362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03355 5361 5362 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03354 7514 5423 5360 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03353 5356 5359 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03352 7514 5356 5336 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03351 5355 5361 5356 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03350 7495 5355 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03349 7514 5355 7495 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03348 5336 5361 5359 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03347 5359 5362 5337 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03346 5623 6344 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03345 7111 1115 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03344 822 1768 821 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03343 820 902 822 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03342 821 1435 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03341 819 822 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03340 7514 899 820 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03339 820 900 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03338 6402 6565 6361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03337 6361 6566 6402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03336 7514 6628 6361 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03335 630 668 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03334 628 670 662 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03333 7514 1168 628 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03332 7514 669 670 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03331 667 670 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03330 7514 841 668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03329 663 665 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03328 7514 663 629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03327 662 667 663 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03326 1168 662 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03325 7514 662 1168 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03324 629 667 665 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03323 665 670 630 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03322 3668 3667 3669 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03321 3669 3743 3668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03320 7514 3836 3669 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03319 3666 3668 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03318 7058 7093 7092 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03317 7514 7094 7058 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03316 7059 7095 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03315 7092 7090 7059 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03314 7514 7095 7093 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03313 7090 7094 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03312 2721 4368 2720 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03311 2720 2733 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03310 2722 4367 2721 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03309 2718 2719 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03308 2719 4724 2722 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03307 4441 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03306 7514 4158 4441 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03305 6992 6491 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03304 5435 5833 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03303 7514 5377 3167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03302 3167 5541 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03301 7514 5378 3167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03300 6656 6679 6678 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03299 7514 6676 6656 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03298 6657 6819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03297 6678 6677 6657 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03296 7514 6819 6679 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03295 6677 6676 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03294 4377 4934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03293 7514 3820 4377 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03292 4592 5842 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03291 4985 7108 4592 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03290 348 370 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03289 7514 953 348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03288 348 372 640 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03287 640 1466 348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03286 3638 3636 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03285 4217 3637 3638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03284 5921 5952 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03283 5954 5953 5921 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03282 5136 5134 5135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03281 5135 5369 5136 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03280 7514 5226 5135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03279 5282 5136 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03278 7514 2934 2714 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03277 2714 5128 2716 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03276 7514 5128 2717 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03275 2716 2717 2715 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03274 2938 2716 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03273 2715 3649 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03272 7514 5075 5029 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03271 5029 5074 5076 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03270 5600 5076 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03269 1107 1211 1108 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03268 1108 4597 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03267 1105 5619 1107 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03266 1106 1709 1105 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03265 2851 3083 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03264 5885 3084 2851 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03263 7514 5125 5126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03262 5126 5128 5129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03261 7514 5128 5131 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03260 5129 5131 5130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03259 5124 5129 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03258 5130 5127 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03257 7514 3475 3477 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03256 3477 5128 3479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03255 7514 5128 3480 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03254 3479 3480 3478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03253 3476 3479 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03252 3478 3804 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03251 7514 3879 3490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03250 3490 5128 3492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03249 7514 5128 3493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03248 3492 3493 3491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03247 3884 3492 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03246 3491 4211 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03245 3321 3501 3320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03244 3320 4669 3321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03243 7514 3644 3320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03242 2038 2814 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03241 2037 2103 2038 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03240 1330 1333 1331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03239 1331 1334 1330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03238 7514 1332 1331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03237 1552 1330 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03236 3031 3033 3034 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03235 3034 3037 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03234 3032 3029 3031 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03233 3738 3030 3032 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03232 4997 4996 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03231 7514 5376 4997 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03230 4997 5087 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03229 7514 4995 4997 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03228 5819 4997 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03227 5133 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03226 5214 7286 5133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03225 5132 5137 5214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03224 7514 5275 5132 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03223 5132 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03222 4302 4448 4301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03221 4301 4441 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03220 4300 4442 4302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03219 5620 4934 4300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03218 1644 2926 1692 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03217 1692 3135 1645 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03216 1645 3012 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03215 1643 2925 1692 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03214 7514 4979 1643 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03213 7514 6173 1644 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03212 1876 1692 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03211 152 183 276 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03210 7514 378 152 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03209 153 771 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03208 276 184 153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03207 7514 771 183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03206 184 378 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03205 5331 5329 5330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03204 5330 6058 5331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03203 7514 5626 5330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03202 4029 6133 4031 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03201 4031 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03200 4030 4158 4029 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03199 4084 4085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03198 4085 7114 4030 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03197 1352 1430 1351 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03196 1351 1723 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03195 1353 1466 1352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03194 2587 1350 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03193 1350 2995 1353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03192 5277 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03191 5411 7286 5277 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03190 5276 5274 5411 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03189 7514 5275 5276 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03188 5276 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03187 538 609 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03186 7514 495 538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03185 538 847 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03184 7514 494 538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03183 1841 538 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03182 5299 5376 5155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03181 5155 5273 5299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03180 7514 5887 5155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03179 6242 6168 6170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03178 6170 6169 6242 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03177 7514 6315 6170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03176 6748 6751 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03175 6744 6753 6745 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03174 7514 7489 6744 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03173 7514 7215 6753 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03172 6752 6753 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03171 7514 6750 6751 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03170 6746 6749 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03169 7514 6746 6747 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03168 6745 6752 6746 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03167 7489 6745 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03166 7514 6745 7489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03165 6747 6752 6749 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03164 6749 6753 6748 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03163 2210 4446 2211 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03162 2211 2880 2268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03161 7514 2881 2210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03160 2687 2268 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03159 6502 6560 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03158 6500 6557 6555 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03157 7514 7466 6500 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03156 7514 6528 6557 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03155 6556 6557 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03154 7514 6561 6560 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03153 6558 6559 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03152 7514 6558 6501 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03151 6555 6556 6558 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03150 7466 6555 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03149 7514 6555 7466 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03148 6501 6556 6559 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03147 6559 6557 6502 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03146 4749 4846 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03145 4765 4764 4749 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03144 4430 4581 4429 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03143 4428 4986 4430 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03142 4429 4427 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03141 4720 4430 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03140 7514 4987 4428 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03139 4428 4984 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_03138 4616 5137 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03137 4920 5832 4616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03136 7514 4649 4920 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03135 7514 6600 6179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03134 7514 6406 6179 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03133 6179 6599 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03132 6180 6179 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03131 5419 5418 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03130 5417 6096 5419 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03129 814 1728 815 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03128 815 937 814 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03127 7514 1681 815 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03126 1333 814 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03125 5237 5207 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03124 7514 5818 5237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03123 5237 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03122 7514 5815 5237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03121 5238 5237 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03120 3191 3411 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03119 4574 3412 3191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03118 5227 5225 5193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03117 5193 5369 5227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03116 7514 5226 5193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03115 5806 5227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03114 4722 4718 4719 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03113 4719 5381 4722 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03112 7514 6386 4719 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03111 2760 2847 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03110 2794 2846 2760 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03109 1910 1915 1909 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03108 1909 1908 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03107 1907 1906 1910 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03106 2748 2686 1907 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03105 5748 5746 5747 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03104 5747 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03103 5749 7042 5748 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03102 6568 7114 5749 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03101 7514 6894 3193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03100 3193 3216 3217 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03099 3304 3217 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03098 7514 606 1051 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03097 606 4934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03096 1051 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03095 7203 7491 7178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03094 7178 7379 7203 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03093 7514 7475 7178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03092 7419 7203 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03091 1357 1355 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03090 1872 1356 1357 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03089 1354 2502 1872 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03088 7514 2435 1354 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03087 1354 2853 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_03086 7514 1444 1383 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03085 7514 1627 1383 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03084 1383 1508 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03083 1382 1383 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03082 7514 4371 4372 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03081 4371 4514 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03080 4372 6600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03079 2984 3633 2985 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03078 2985 2999 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03077 2983 3632 2984 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03076 3216 2998 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03075 2998 3300 2983 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03074 7514 6333 5346 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03073 5346 5457 5382 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03072 6979 5382 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03071 2196 2418 2197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03070 2197 2222 2223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03069 7514 2220 2196 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03068 2221 2223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_03067 2442 2664 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03066 3005 5882 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03065 1346 1349 1550 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03064 7514 1427 1346 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03063 1348 1558 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03062 1550 1347 1348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03061 7514 1558 1349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03060 1347 1427 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03059 3964 4437 3965 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03058 3965 4081 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03057 3963 6266 3964 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03056 4511 3999 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_03055 3999 7162 3963 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03054 5173 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03053 7514 2111 5173 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03052 5207 5160 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03051 2517 2934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03050 4838 5137 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03049 2165 3418 2166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03048 2166 2929 2165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03047 7514 5882 2166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03046 3781 3783 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03045 3775 3784 3776 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03044 7514 3774 3775 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03043 7514 4638 3784 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03042 3782 3784 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_03041 7514 3779 3783 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_03040 3777 3780 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03039 7514 3777 3778 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03038 3776 3782 3777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03037 3774 3776 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03036 7514 3776 3774 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03035 3778 3782 3780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03034 3780 3784 3781 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03033 2574 2688 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03032 2825 2687 2574 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03031 7514 4627 4629 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03030 4627 4833 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03029 4629 4752 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03028 7395 7415 7416 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03027 7514 7465 7395 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03026 7394 7418 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03025 7416 7414 7394 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03024 7514 7418 7415 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03023 7414 7465 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_03022 1249 1577 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03021 1287 5000 1249 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03020 5474 5505 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03019 5723 5506 5474 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03018 2627 2659 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03017 3084 2707 2627 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03016 7514 3086 2765 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03015 2765 4106 2805 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03014 7514 4106 2807 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03013 2805 2807 2766 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03012 3092 2805 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03011 2766 3649 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03010 7514 4104 4105 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03009 4105 4106 4108 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03008 7514 4106 4109 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03007 4108 4109 4107 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03006 4103 4108 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_03005 4107 5127 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03004 1897 2814 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03003 1896 2811 1897 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_03002 7514 3696 3672 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03001 3672 4106 3698 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_03000 7514 4106 3700 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02999 3698 3700 3673 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02998 3695 3698 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02997 3673 3804 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02996 7514 4113 3675 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02995 3675 4106 3708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02994 7514 4106 3709 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02993 3708 3709 3676 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02992 4119 3708 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02991 3676 4211 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02990 7514 4921 4879 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02989 4879 4920 4922 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02988 5521 4922 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02987 5612 5969 5613 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02986 5613 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02985 5611 5841 5612 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02984 6399 7114 5611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02983 5544 7390 5492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02982 7514 7388 5545 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02981 5492 5545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02980 2780 5994 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02979 2823 6133 2780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02978 2779 6266 2823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02977 7514 5840 2779 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02976 2779 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02975 7067 7431 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02974 7123 7107 7067 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02973 834 960 835 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02972 835 832 834 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02971 7514 2592 835 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02970 833 834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02969 1260 1732 1221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02968 1221 1547 1260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02967 7514 1548 1221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02966 2007 1260 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02965 3131 3129 3130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02964 3130 4695 3131 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02963 7514 3128 3130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02962 6042 6565 6043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02961 6043 6566 6042 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02960 7514 6676 6043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02959 6471 7227 6470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02958 6470 7228 6471 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02957 7514 7466 6470 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02956 6088 6843 6089 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02955 6089 6405 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02954 6087 6768 6088 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02953 7034 6132 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02952 6132 6907 6087 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02951 6094 6372 6067 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02950 6067 6293 6094 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02949 7514 7420 6067 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02948 6185 7227 6186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02947 6186 7228 6185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02946 7514 7493 6186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02945 6866 6867 7011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02944 7514 7453 6866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02943 6868 7074 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02942 7011 6865 6868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02941 7514 7074 6867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02940 6865 7453 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02939 37 39 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02938 32 40 33 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02937 7514 6266 32 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02936 7514 403 40 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02935 38 40 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02934 7514 41 39 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02933 34 36 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02932 7514 34 35 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02931 33 38 34 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02930 6266 33 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02929 7514 33 6266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02928 35 38 36 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02927 36 40 37 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02926 7514 5889 5037 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02925 5037 5844 5094 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02924 5093 5094 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02923 7514 2182 2184 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02922 2184 2183 2186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02921 2185 2186 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02920 7514 1976 1905 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02919 1905 4448 1904 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02918 2322 1904 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02917 3816 3890 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02916 7105 4228 3816 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02915 3815 3814 7105 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02914 7514 4149 3815 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02913 3815 5909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02912 2508 3418 2296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02911 2296 2929 2508 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02910 7514 6025 2296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02909 2075 2383 2076 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02908 2076 2514 2096 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02907 7514 2304 2075 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02906 2095 2096 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02905 4157 4156 4159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02904 7514 4158 4160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02903 4159 4160 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02902 7514 7384 5910 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02901 5910 7286 5911 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02900 5909 5911 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02899 6731 7280 6730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02898 6730 7428 6731 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02897 7514 6965 6730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02896 970 972 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02895 965 973 964 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02894 7514 963 965 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02893 7514 1290 973 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02892 971 973 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02891 7514 968 972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02890 966 969 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02889 7514 966 967 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02888 964 971 966 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02887 963 964 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02886 7514 964 963 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02885 967 971 969 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02884 969 973 970 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02883 3732 3742 3376 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02882 3376 3425 3732 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02881 7514 4148 3376 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02880 6593 6166 6167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02879 6167 6165 6593 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02878 7514 6315 6167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02877 1935 4568 1936 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02876 1936 2452 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02875 1934 4588 1935 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02874 1968 1969 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02873 1969 4569 1934 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02872 2684 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02871 7514 4161 2684 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02870 1167 2543 1140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02869 1140 2541 1167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02868 7514 1445 1140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02867 1837 1167 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02866 4166 4173 4167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02865 4165 4175 4166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02864 4937 4166 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02863 7514 4166 4937 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02862 4171 4174 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02861 7514 4172 4174 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02860 4173 4175 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02859 7514 4305 4175 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02858 4168 4170 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02857 4167 7500 4168 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02856 4170 4175 4171 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02855 4169 4173 4170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02854 7514 4167 4169 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02853 7514 4937 4164 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02852 4164 7500 4165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02851 4750 5072 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02850 4774 4773 4750 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02849 5940 6133 5941 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02848 5941 5994 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02847 6843 7114 5940 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02846 6968 6599 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02845 7514 6848 6968 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02844 6968 6600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02843 7514 6981 6968 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02842 4970 4971 4972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02841 4972 5369 4970 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02840 7514 5226 4972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02839 5801 4970 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02838 2626 3213 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02837 2658 2657 2626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02836 1442 1441 1409 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02835 1409 1440 1442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02834 7514 4597 1409 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02833 1759 1442 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02832 845 1908 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02831 844 1915 845 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02830 3425 2686 2572 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02829 7514 4934 2611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02828 2572 2611 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02827 3812 3811 3813 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02826 3813 4360 3812 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02825 7514 6041 3813 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02824 3810 3812 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02823 6024 6968 6022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02822 6022 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02821 6023 7462 6024 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02820 7152 7280 7153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02819 7153 7428 7152 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02818 7514 7493 7153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02817 7151 7152 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02816 2204 2255 2205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02815 2205 2390 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02814 2608 7162 2204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02813 7514 4588 4188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02812 4188 4297 4230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02811 4231 4230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02810 1082 2842 1081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02809 1081 2792 1082 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02808 7514 2133 1081 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02807 2155 2154 2156 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02806 2156 2434 2155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02805 7514 2164 2156 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02804 2153 2155 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02803 3060 4437 3059 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02802 3059 4600 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02801 3058 6133 3060 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02800 4588 7114 3058 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02799 6792 7164 6793 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02798 6793 6914 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02797 6791 7286 6792 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02796 6839 7113 6791 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02795 5031 6832 5032 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02794 5032 5079 5080 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02793 7514 5238 5031 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02792 5078 5080 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02791 1659 1915 1660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02790 1660 1908 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02789 1658 1906 1659 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02788 1767 4000 1658 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02787 1233 4081 1232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02786 1232 1292 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02785 1231 5001 1233 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02784 4569 5690 1231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02783 7514 5996 7384 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02782 5996 6652 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02781 7384 6061 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02780 2055 4694 2056 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02779 2056 2141 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02778 2054 2524 2055 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02777 2085 2228 2054 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02776 6049 6048 6051 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02775 6051 6193 6050 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02774 7514 6046 6049 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02773 6047 6050 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02772 7166 7391 7165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02771 7165 7164 7167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02770 7514 7162 7166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02769 7163 7167 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02768 6066 6118 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02767 6064 6121 6115 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02766 7514 7452 6064 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02765 7514 6231 6121 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02764 6120 6121 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02763 7514 6119 6118 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02762 6116 6117 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02761 7514 6116 6065 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02760 6115 6120 6116 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02759 7452 6115 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02758 7514 6115 7452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02757 6065 6120 6117 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02756 6117 6121 6066 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02755 4649 4502 4461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02754 4461 5381 4649 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02753 7514 6386 4461 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02752 2703 3149 2704 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02751 2704 4695 2703 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02750 7514 3213 2704 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02749 2847 2703 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02748 7514 3167 472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02747 434 472 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02746 7514 472 434 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02745 7514 472 434 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02744 434 472 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02743 7514 434 386 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02742 1688 386 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02741 7514 386 1688 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02740 7514 386 1688 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02739 1688 386 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02738 7514 434 328 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02737 3546 328 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02736 7514 328 3546 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02735 7514 328 3546 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02734 3546 328 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02733 7514 579 285 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02732 331 285 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02731 7514 285 331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02730 7514 285 331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02729 331 285 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02728 7514 331 332 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02727 3352 332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02726 7514 332 3352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02725 7514 332 3352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02724 3352 332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02723 7514 331 228 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02722 4934 228 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02721 7514 228 4934 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02720 7514 228 4934 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02719 4934 228 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02718 5873 5872 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02717 5867 5874 5866 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02716 7514 6628 5867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02715 7514 6302 5874 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02714 5875 5874 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02713 7514 5870 5872 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02712 5868 5871 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02711 7514 5868 5869 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02710 5866 5875 5868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02709 6628 5866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02708 7514 5866 6628 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02707 5869 5875 5871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02706 5871 5874 5873 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02705 2339 2337 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02704 7514 2338 2339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02703 2339 2467 2456 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02702 2456 3837 2339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02701 6494 6543 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02700 6492 6545 6540 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02699 7514 6539 6492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02698 7514 6622 6545 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02697 6544 6545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02696 7514 6549 6543 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02695 6546 6542 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02694 7514 6546 6493 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02693 6540 6544 6546 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02692 6539 6540 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02691 7514 6540 6539 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02690 6493 6544 6542 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02689 6542 6545 6494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02688 7514 2167 4697 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02687 2167 2168 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02686 4697 3214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02685 4696 4104 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02684 5134 4834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02683 3771 6432 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02682 7514 6714 6538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02681 6538 6852 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02680 7514 7113 6538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02679 1198 1287 1199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02678 1199 1823 1198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02677 7514 1197 1199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02676 2029 1198 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02675 2448 2449 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02674 2443 2451 2444 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02673 7514 2602 2443 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02672 7514 2533 2451 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02671 2450 2451 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02670 7514 2603 2449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02669 2445 2446 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02668 7514 2445 2447 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02667 2444 2450 2445 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02666 2602 2444 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02665 7514 2444 2602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02664 2447 2450 2446 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02663 2446 2451 2448 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02662 5653 5969 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02661 4112 6175 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02660 5175 5171 5176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02659 5176 5172 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02658 5174 5173 5175 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02657 5457 5170 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02656 5170 6266 5174 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02655 7514 4411 3846 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02654 3846 4197 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02653 3878 3877 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02652 3846 4413 3877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02651 3877 4908 3846 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02650 2392 4158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02649 7514 3352 2392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02648 354 4517 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02647 495 405 354 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02646 1730 3979 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02645 1728 1727 1730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02644 1729 3546 1728 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02643 7514 2139 1729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02642 1729 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02641 5771 5809 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02640 5960 5877 5771 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02639 7078 7280 7054 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02638 7054 7428 7078 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02637 7514 7453 7054 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02636 7514 4504 3367 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02635 3367 4264 3417 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02634 7514 4264 3388 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02633 3417 3388 3366 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02632 3582 3417 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02631 3366 3387 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02630 1218 3469 1217 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02629 1217 3472 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02628 5127 3470 1218 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02627 7514 4502 3150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02626 3150 4264 3151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02625 7514 4264 3153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02624 3151 3153 3152 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02623 3315 3151 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02622 3152 3410 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02621 7514 4716 4262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02620 4262 4264 4263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02619 7514 4264 4267 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02618 4263 4267 4266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02617 4261 4263 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02616 4266 4265 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02615 950 1700 952 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02614 952 1968 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02613 951 1435 950 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02612 4830 4828 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02611 4829 6266 4830 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02610 2148 2507 2147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02609 2147 3769 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02608 2416 2508 2148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02607 7514 3347 2876 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02606 2876 4372 2877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02605 2875 2877 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02604 7514 4861 3494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02603 3494 4264 3497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02602 7514 4264 3498 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02601 3497 3498 3496 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02600 3797 3497 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02599 3496 3495 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_02598 1815 1869 1786 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02597 1785 3546 1815 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02596 1786 3000 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02595 1813 1815 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02594 7514 2095 1785 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02593 1785 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02592 3691 5173 3692 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02591 3692 5172 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02590 3690 4446 3691 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02589 3744 3742 3690 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02588 5636 5660 5637 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02587 5637 6094 5661 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02586 7514 5803 5636 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02585 5659 5661 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02584 2948 2945 2901 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02583 2901 2946 2948 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02582 7514 5055 2901 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02581 6189 6187 6190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02580 6190 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02579 6188 7042 6189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02578 6572 6333 6188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02577 7514 7114 1011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02576 1011 1837 1045 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02575 1044 1045 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02574 7514 6181 5934 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02573 5934 5985 5986 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02572 5984 5986 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02571 1927 3012 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02570 2159 3135 1927 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02569 1926 2926 2159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02568 7514 6173 1926 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02567 1925 2925 2159 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02566 7514 4979 1925 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02565 5779 6328 5780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02564 5780 5835 5836 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02563 7514 6471 5779 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02562 5834 5836 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02561 1189 2842 1188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02560 1188 2792 1189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02559 7514 2133 1188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02558 1187 1189 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02557 7514 7114 1656 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02556 1656 1833 1706 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02555 2035 1706 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02554 6796 6980 6797 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02553 6797 6979 6842 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02552 7514 7480 6796 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02551 6841 6842 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02550 6666 6764 6667 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02549 6667 6705 6706 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02548 7514 6899 6666 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02547 6704 6706 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02546 5503 6166 5272 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02545 5272 6165 5503 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02544 7514 5876 5272 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02543 6663 6691 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02542 6661 6694 6685 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02541 7514 7494 6661 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02540 7514 6693 6694 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02539 6695 6694 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02538 7514 6690 6691 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02537 6687 6688 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02536 7514 6687 6662 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02535 6685 6695 6687 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02534 7494 6685 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02533 7514 6685 7494 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02532 6662 6695 6688 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02531 6688 6694 6663 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02530 7370 7368 7372 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02529 7514 7369 7370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02528 7373 7477 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02527 7372 7371 7373 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02526 7514 7477 7368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02525 7371 7369 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02524 5738 6168 5737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02523 5737 6169 5738 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02522 7514 5815 5737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02521 1135 1775 1136 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02520 1136 5171 1165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02519 7514 2881 1135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02518 1501 1165 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02517 4791 5842 4747 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02516 4747 5691 4791 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02515 7514 6133 4747 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02514 4790 4791 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02513 2848 2846 2849 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02512 2849 2991 2850 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02511 2850 2995 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02510 2845 2931 2849 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02509 7514 4254 2845 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02508 7514 2847 2848 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02507 2844 2849 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02506 992 1027 1146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02505 7514 1732 992 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02504 993 1149 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02503 1146 1026 993 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02502 7514 1149 1027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02501 1026 1732 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02500 6926 6975 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02499 6924 6974 6971 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02498 7514 7480 6924 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02497 7514 7225 6974 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02496 6977 6974 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02495 7514 6976 6975 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02494 6972 6973 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02493 7514 6972 6925 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02492 6971 6977 6972 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02491 7480 6971 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02490 7514 6971 7480 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02489 6925 6977 6973 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02488 6973 6974 6926 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02487 5201 5230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02486 5229 5366 5201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02485 2769 3810 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02484 2810 3013 2769 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02483 3036 6133 3035 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02482 3035 5994 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02481 3119 5000 3036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02480 570 1082 572 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02479 572 771 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02478 571 3546 570 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02477 1532 2033 1533 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02476 1533 1570 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02475 1531 4600 1532 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02474 2102 5690 1531 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02473 5755 6048 5754 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02472 5754 6193 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02471 6599 6046 5755 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02470 3021 4437 3022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02469 3022 4081 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02468 3020 6266 3021 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02467 4773 7162 3020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02466 217 220 372 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02465 7514 276 217 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02464 219 280 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02463 372 218 219 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02462 7514 280 220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02461 218 276 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02460 5770 5806 5769 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02459 5769 6162 5808 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02458 7514 5807 5770 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02457 5805 5808 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02456 1752 1880 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02455 2865 1876 1752 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02454 1751 1749 2865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02453 7514 1750 1751 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02452 1748 1746 2865 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02451 7514 1747 1748 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02450 6834 7033 6787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02449 6788 6886 6834 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02448 6787 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02447 6832 6834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02446 7514 7032 6788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02445 6788 7313 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02444 5647 6266 5646 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02443 5646 6332 5689 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02442 7514 7114 5647 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02441 5688 5689 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02440 7514 5897 5308 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02439 5308 5306 5309 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02438 5307 5309 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02437 7514 3637 3365 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02436 3365 3636 3414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02435 3495 3414 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02434 7514 3406 3363 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02433 3363 3407 3408 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02432 3562 3408 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02431 7514 1577 1130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02430 1130 2816 1160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02429 1159 1160 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02428 5421 5735 5027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02427 5027 5734 5421 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02426 7514 5069 5027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02425 7514 4589 4286 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02424 4286 4588 4287 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02423 4583 4287 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02422 7514 1435 1089 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02421 1089 1768 1088 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02420 1466 1088 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02419 551 2290 553 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02418 552 3546 551 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02417 553 3625 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02416 1636 551 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02415 7514 3549 552 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02414 552 1866 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02413 7514 3322 3197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02412 3197 4066 3234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02411 3233 3234 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02410 7514 7042 6800 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02409 6800 7109 6844 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02408 7334 6844 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02407 7514 1775 985 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02406 985 5171 986 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02405 4437 986 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02404 2143 3023 2144 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02403 2142 2292 2143 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02402 2144 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02401 2140 2143 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02400 7514 2141 2142 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02399 2142 2139 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_02398 956 1968 957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02397 957 2718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02396 955 1700 956 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02395 953 954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02394 954 1688 955 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02393 4971 5274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02392 3129 3868 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02391 3149 3774 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02390 4841 5055 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02389 3481 3696 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02388 61 4437 62 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02387 62 4081 111 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02386 7514 6266 61 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02385 195 111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02384 1184 1548 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02383 1182 1952 1184 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02382 1183 1337 1182 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02381 7514 1419 1183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02380 1183 1336 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02379 4330 4377 4331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02378 4331 4447 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02377 4329 4442 4330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02376 7109 4374 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02375 4374 4376 4329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02374 3070 2288 2289 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02373 2289 2287 3070 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02372 7514 2784 2289 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02371 6615 6614 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02370 6613 6851 6615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02369 5914 5912 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02368 5913 7162 5914 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02367 5953 6316 5473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02366 5473 6314 5953 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02365 7514 5876 5473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02364 6649 7286 6650 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02363 6650 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02362 6648 7496 6649 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02361 5675 5884 5342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02360 5342 5885 5675 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02359 7514 5815 5342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02358 996 1035 5884 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02357 7514 1032 996 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02356 995 1034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02355 5884 1031 995 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02354 7514 1034 1035 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02353 1031 1032 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02352 3013 3501 3014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02351 3014 4669 3013 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02350 7514 3012 3014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02349 1930 4588 1929 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02348 1929 4568 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02347 2926 4569 1930 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02346 7514 988 1915 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02345 988 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02344 1915 2111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02343 6367 6906 6368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02342 6368 6710 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02341 6366 6407 6367 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02340 6409 6408 6366 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02339 3649 4987 3330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02338 3330 4984 3649 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02337 7514 4986 3330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02336 7142 7280 7143 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02335 7143 7428 7142 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02334 7514 7466 7143 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02333 7210 7142 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02332 3576 3583 3577 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02331 3532 3585 3576 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02330 4504 3576 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02329 7514 3576 4504 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02328 3534 3584 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02327 7514 3582 3584 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02326 3583 3585 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02325 7514 3581 3585 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02324 3531 3579 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02323 3577 7500 3531 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02322 3579 3585 3534 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02321 3533 3583 3579 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02320 7514 3577 3533 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02319 7514 4504 3530 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02318 3530 7500 3532 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02317 4738 5216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02316 5074 5832 4738 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02315 7514 4769 5074 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02314 7514 1694 1490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02313 1490 1489 1491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02312 3160 1491 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02311 7514 7286 6330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02310 6330 7164 6331 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02309 6981 6331 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02308 7514 4665 4780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02307 4665 4726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02306 4780 4995 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02305 7514 4367 4319 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02304 4319 4368 4369 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02303 4781 4369 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02302 7514 4569 3373 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02301 3373 4568 3421 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02300 3420 3421 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02299 7514 6324 6326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02298 6324 6325 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02297 6326 6757 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02296 1197 2435 1126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02295 1126 2853 1197 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02294 7514 2504 1126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02293 6218 7042 6219 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02292 6219 6332 6265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02291 7514 7162 6218 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02290 6338 6265 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02289 2900 2942 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02288 2898 2944 2936 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02287 7514 2934 2898 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02286 7514 3571 2944 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02285 2943 2944 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02284 7514 2938 2942 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02283 2937 2940 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02282 7514 2937 2899 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02281 2936 2943 2937 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02280 2934 2936 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02279 7514 2936 2934 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02278 2899 2943 2940 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02277 2940 2944 2900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02276 5099 5106 5101 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02275 5039 5107 5099 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02274 7388 5099 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02273 7514 5099 7388 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02272 5042 5105 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02271 7514 5393 5105 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02270 5106 5107 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02269 7514 5554 5107 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02268 5040 5103 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02267 5101 5100 5040 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02266 5103 5107 5042 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02265 5041 5106 5103 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02264 7514 5101 5041 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02263 7514 7388 5038 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02262 5038 5100 5039 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02261 5352 6316 4875 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02260 4875 6314 5352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02259 7514 5069 4875 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02258 5710 5711 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02257 5974 5738 5710 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02256 5789 6061 5788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02255 5788 6652 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02254 5787 7390 5789 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02253 5912 5845 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_02252 5845 7388 5787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02251 1420 1333 1335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02250 1335 1334 1420 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02249 7514 1332 1335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02248 2004 2005 5735 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02247 7514 2002 2004 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02246 2006 2082 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02245 5735 2003 2006 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02244 7514 2082 2005 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02243 2003 2002 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02242 3736 3922 3378 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02241 3378 3925 3736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02240 7514 5055 3378 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02239 2180 2543 2181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02238 2181 2541 2180 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02237 7514 2179 2181 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02236 2390 2180 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02235 7514 2221 3472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02234 3472 2366 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02233 7514 2217 3472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02232 6955 7227 6927 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02231 6927 7228 6955 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02230 7514 7464 6927 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02229 4721 5078 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02228 4857 4720 4721 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02227 6077 6992 6078 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02226 6078 6410 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02225 6202 6135 6077 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02224 6124 7491 5925 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02223 5925 7379 6124 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02222 7514 6676 5925 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02221 6306 6393 6174 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02220 6174 6394 6306 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02219 7514 6173 6174 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02218 6755 6968 6754 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02217 6754 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02216 6837 7480 6755 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02215 2855 3135 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02214 2854 3645 2855 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02213 7514 5695 5469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02212 5469 5544 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02211 6056 5468 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02210 5469 5466 5468 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02209 5468 5467 5469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_02208 448 3346 447 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02207 447 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02206 446 1304 448 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02205 240 3346 241 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02204 241 2887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02203 239 1906 240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02202 5487 5536 5486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02201 5486 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02200 5485 5841 5487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02199 5985 7162 5485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02198 2710 3710 2711 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02197 2711 4695 2710 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02196 7514 3145 2711 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02195 2800 2710 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02194 3654 3656 4074 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02193 7514 5138 3654 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02192 3657 3655 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02191 4074 3653 3657 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02190 7514 3655 3656 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02189 3653 5138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02188 7060 7493 7061 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02187 7061 7489 7096 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02186 7514 7494 7060 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02185 7095 7096 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02184 5813 6166 5773 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02183 5773 6165 5813 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02182 7514 5815 5773 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02181 2521 2945 2441 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02180 2441 2946 2521 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02179 7514 4834 2441 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02178 1547 1146 818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02177 818 1182 1547 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02176 7514 1145 818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02175 6380 7491 6350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02174 6350 7379 6380 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02173 7514 6628 6350 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02172 5722 5724 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02171 5704 5726 5721 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02170 7514 7454 5704 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02169 7514 6231 5726 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02168 5725 5726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02167 7514 5723 5724 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02166 5705 5706 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02165 7514 5705 5707 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02164 5721 5725 5705 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02163 7454 5721 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02162 7514 5721 7454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02161 5707 5725 5706 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02160 5706 5726 5722 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02159 7514 951 946 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02158 946 949 947 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02157 1145 947 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02156 7514 6402 6074 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02155 6074 6128 6129 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02154 6325 6129 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02153 1913 1914 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02152 2325 1911 1913 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02151 1912 2536 2325 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02150 7514 2398 1912 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02149 1912 2813 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02148 7514 2602 2203 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02147 2203 4161 2251 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02146 2811 2251 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02145 7016 7491 7017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02144 7017 7379 7016 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02143 7514 7462 7017 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02142 5762 5798 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02141 5760 5800 5792 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02140 7514 6965 5760 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02139 7514 6231 5800 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02138 5799 5800 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02137 7514 5797 5798 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02136 5793 5794 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02135 7514 5793 5761 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02134 5792 5799 5793 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02133 6965 5792 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02132 7514 5792 6965 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02131 5761 5799 5794 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02130 5794 5800 5762 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02129 1192 1700 1191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02128 1191 1968 1226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02127 7514 1435 1192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02126 1866 1226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_02125 6205 6228 6226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02124 7514 7335 6205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02123 6206 6726 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02122 6226 6225 6206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02121 7514 6726 6228 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02120 6225 7335 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02119 4965 4968 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02118 4960 4969 4961 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02117 7514 4959 4960 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02116 7514 5584 4969 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02115 4967 4969 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02114 7514 4966 4968 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_02113 4962 4963 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02112 7514 4962 4964 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02111 4961 4967 4962 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02110 4959 4961 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02109 7514 4961 4959 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02108 4964 4967 4963 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02107 4963 4969 4965 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02106 4151 4207 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02105 5989 4228 4151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02104 4150 4148 5989 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02103 7514 4149 4150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02102 4150 5909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_02101 1440 1906 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02100 7514 1304 1440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_02099 7465 7464 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02098 4412 6035 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02097 5371 5536 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02096 7514 3210 3133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02095 3132 3133 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02094 7514 3133 3132 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02093 7514 3133 3132 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02092 3132 3133 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02091 7514 3210 3205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02090 3204 3205 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02089 7514 3205 3204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02088 7514 3205 3204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02087 3204 3205 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02086 7514 3210 3206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02085 3400 3206 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02084 7514 3206 3400 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02083 7514 3206 3400 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02082 3400 3206 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02081 7514 3210 3141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02080 3140 3141 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02079 7514 3141 3140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02078 7514 3141 3140 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02077 3140 3141 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02076 7514 3210 3209 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02075 3208 3209 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02074 7514 3209 3208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02073 7514 3209 3208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02072 3208 3209 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02071 7514 3210 3211 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02070 3558 3211 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02069 7514 3211 3558 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02068 7514 3211 3558 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02067 3558 3211 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02066 7514 3229 2152 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02065 2151 2152 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02064 7514 2152 2151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02063 7514 2152 2151 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02062 2151 2152 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02061 2698 2926 2700 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02060 2700 3135 2699 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02059 2699 3644 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02058 2697 2925 2700 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02057 7514 5216 2697 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02056 7514 6388 2698 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02055 2696 2700 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02054 6733 6676 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02053 3811 3727 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02052 5204 5616 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02051 5837 5457 5204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02050 6211 6309 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02049 6561 6246 6211 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02048 7514 3229 2233 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02047 2232 2233 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02046 7514 2233 2232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02045 7514 2233 2232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02044 2232 2233 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02043 7514 3229 2235 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02042 2234 2235 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02041 7514 2235 2234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02040 7514 2235 2234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02039 2234 2235 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02038 7514 3229 2162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02037 2163 2162 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02036 7514 2162 2163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02035 7514 2162 2163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02034 2163 2162 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02033 7514 3229 2238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02032 2237 2238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02031 7514 2238 2237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02030 7514 2238 2237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02029 2237 2238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02028 7514 3229 2240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02027 2239 2240 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02026 7514 2240 2239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02025 7514 2240 2239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02024 2239 2240 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02023 7514 3229 3148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02022 3147 3148 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02021 7514 3148 3147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02020 7514 3148 3147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02019 3147 3148 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02018 7514 3229 3219 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02017 3218 3219 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02016 7514 3219 3218 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02015 7514 3219 3218 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02014 3218 3219 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02013 7514 3229 3221 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02012 3220 3221 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02011 7514 3221 3220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02010 7514 3221 3220 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02009 3220 3221 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02008 7275 7277 7274 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02007 7514 7480 7275 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02006 7276 7477 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02005 7274 7273 7276 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_02004 7514 7477 7277 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02003 7273 7480 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_02002 2497 2785 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02001 2505 2837 2497 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_02000 7514 6852 6715 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01999 6715 6714 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01998 6849 6715 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01997 5823 5817 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01996 7514 5818 5823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01995 5823 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01994 7514 5815 5823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01993 5816 5823 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01992 5599 6637 5602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01991 5602 5600 5601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01990 7514 5669 5599 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01989 5711 5601 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01988 3203 5691 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01987 3266 5001 3203 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01986 2478 3769 2479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01985 2479 2583 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01984 2477 2507 2478 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01983 2653 2508 2477 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01982 7514 3229 3154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01981 3155 3154 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01980 7514 3154 3155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01979 7514 3154 3155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01978 3155 3154 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01977 7514 3229 3228 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01976 3227 3228 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01975 7514 3228 3227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01974 7514 3228 3227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01973 3227 3228 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01972 7514 3229 3230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01971 3571 3230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01970 7514 3230 3571 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01969 7514 3230 3571 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01968 3571 3230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01967 7514 2712 852 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01966 1264 852 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01965 7514 852 1264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01964 7514 852 1264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01963 1264 852 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01962 1506 1915 1505 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01961 1505 1908 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01960 1835 1906 1506 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01959 7514 1054 4448 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01958 1054 4376 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01957 4448 3820 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01956 6344 7235 5942 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01955 7514 6652 5995 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01954 5942 5995 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01953 210 1025 209 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01952 209 266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01951 1216 1543 210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01950 1689 1876 1665 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01949 1664 1688 1689 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01948 1665 1851 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01947 1686 1689 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01946 7514 2095 1664 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01945 1664 3545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01944 6873 7335 6872 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01943 6872 7074 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01942 6871 7452 6873 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01941 6869 6870 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01940 6870 7453 6871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01939 7514 2712 856 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01938 1281 856 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01937 7514 856 1281 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01936 7514 856 1281 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01935 1281 856 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01934 7514 2712 2701 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01933 3210 2701 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01932 7514 2701 3210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01931 7514 2701 3210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01930 3210 2701 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01929 7514 2712 2713 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01928 3229 2713 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01927 7514 2713 3229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01926 7514 2713 3229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01925 3229 2713 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01924 7149 7151 7150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01923 7150 7315 7149 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01922 7514 7420 7150 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01921 4047 4054 4050 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01920 4011 4053 4047 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01919 4716 4047 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01918 7514 4047 4716 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01917 4014 4052 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01916 7514 4261 4052 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01915 4054 4053 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01914 7514 4488 4053 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01913 4012 4048 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01912 4050 7500 4012 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01911 4048 4053 4014 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01910 4013 4054 4048 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01909 7514 4050 4013 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01908 7514 4716 4010 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01907 4010 7500 4011 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01906 3601 3922 3543 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01905 3543 3925 3601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01904 7514 5274 3543 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01903 7514 1295 330 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01902 329 330 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01901 7514 330 329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01900 7514 330 329 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01899 329 330 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01898 7514 1295 388 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01897 387 388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01896 7514 388 387 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01895 7514 388 387 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01894 387 388 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01893 7514 1295 389 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01892 788 389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01891 7514 389 788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01890 7514 389 788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01889 788 389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01888 7514 1295 334 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01887 333 334 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01886 7514 334 333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01885 7514 334 333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01884 333 334 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01883 7514 1295 393 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01882 392 393 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01881 7514 393 392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01880 7514 393 392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01879 392 393 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01878 7514 1295 394 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01877 598 394 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01876 7514 394 598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01875 7514 394 598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01874 598 394 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01873 7514 1295 1230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01872 1201 1230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01871 7514 1230 1201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01870 7514 1230 1201 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01869 1201 1230 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01868 7514 3719 3681 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01867 3681 4142 3721 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01866 3720 3721 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01865 1162 1368 1132 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01864 1131 1365 1162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01863 1132 4437 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01862 1971 1162 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01861 7514 1366 1131 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01860 1131 1500 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01859 7514 4158 2357 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01858 2357 4934 2389 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01857 2816 2389 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01856 7514 7388 7301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01855 7301 7390 7336 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01854 7353 7336 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01853 7514 1111 873 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01852 873 1109 917 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01851 1620 917 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01850 3213 3214 3192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01849 3192 3212 3213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01848 7514 3550 3192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01847 7514 1295 1289 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01846 1288 1289 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01845 7514 1289 1288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01844 7514 1289 1288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01843 1288 1289 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01842 7514 1295 1291 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01841 1290 1291 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01840 7514 1291 1290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01839 7514 1291 1290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01838 1290 1291 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01837 7514 1295 1234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01836 1206 1234 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01835 7514 1234 1206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01834 7514 1234 1206 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01833 1206 1234 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01832 7514 1295 1293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01831 1294 1293 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01830 7514 1293 1294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01829 7514 1293 1294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01828 1294 1293 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01827 7514 1295 1297 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01826 1296 1297 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01825 7514 1297 1296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01824 7514 1297 1296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01823 1296 1297 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01822 7514 1310 336 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01821 335 336 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01820 7514 336 335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01819 7514 336 335 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01818 335 336 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01817 7514 1310 397 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01816 396 397 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01815 7514 397 396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01814 7514 397 396 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01813 396 397 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01812 7514 1310 398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01811 669 398 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01810 7514 398 669 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01809 7514 398 669 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01808 669 398 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01807 4559 4560 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01806 4554 4563 4555 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01805 7514 6173 4554 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01804 7514 4561 4563 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01803 4562 4563 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01802 7514 4644 4560 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01801 4556 4557 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01800 7514 4556 4558 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01799 4555 4562 4556 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01798 6173 4555 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01797 7514 4555 6173 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01796 4558 4562 4557 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01795 4557 4563 4559 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01794 1008 4600 1009 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01793 1009 1292 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01792 1007 5001 1008 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01791 1569 1042 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01790 1042 5690 1007 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01789 1380 1581 1381 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01788 1381 1631 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01787 1379 1377 1380 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01786 1376 1378 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01785 1378 1618 1379 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01784 492 4600 491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01783 491 1292 532 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01782 7514 6266 492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01781 533 532 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01780 2538 2543 2492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01779 2492 2541 2538 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01778 7514 2542 2492 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01777 2537 2538 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01776 6801 6846 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01775 7514 6845 6801 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01774 6801 6849 6848 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01773 6848 7287 6801 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01772 4892 5171 4893 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01771 4893 5172 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01770 4891 5173 4892 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01769 6565 4936 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01768 4936 6133 4891 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01767 4606 5842 4605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01766 4605 5691 4606 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01765 7514 5841 4605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01764 4604 4606 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01763 7107 6314 6071 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01762 6071 6316 7107 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01761 7514 6125 6071 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01760 7514 1310 344 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01759 343 344 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01758 7514 344 343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01757 7514 344 343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01756 343 344 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01755 7514 1310 402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01754 401 402 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01753 7514 402 401 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01752 7514 402 401 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01751 401 402 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01750 7514 1310 404 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01749 403 404 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01748 7514 404 403 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01747 7514 404 403 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01746 403 404 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01745 7514 1310 1238 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01744 1210 1238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01743 7514 1238 1210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01742 7514 1238 1210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01741 1210 1238 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01740 7514 1310 1301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01739 1300 1301 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01738 7514 1301 1300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01737 7514 1301 1300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01736 1300 1301 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01735 7514 1310 1303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01734 1302 1303 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01733 7514 1303 1302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01732 7514 1303 1302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01731 1302 1303 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01730 7514 1310 1244 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01729 1215 1244 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01728 7514 1244 1215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01727 7514 1244 1215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01726 1215 1244 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01725 4769 4716 4717 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01724 4717 5381 4769 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01723 7514 6386 4717 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01722 1527 1568 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01721 2168 1569 1527 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01720 5012 4589 4025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01719 4025 4074 5012 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01718 7514 4075 4025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01717 4840 4838 4839 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01716 4839 5369 4840 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01715 7514 5226 4839 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01714 5728 4840 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01713 7436 7443 7437 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01712 7405 7444 7436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01711 7512 7436 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01710 7514 7436 7512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01709 7408 7442 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01708 7514 7440 7442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01707 7443 7444 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01706 7514 7508 7444 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01705 7406 7439 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01704 7437 7500 7406 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01703 7439 7444 7408 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01702 7407 7443 7439 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01701 7514 7437 7407 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01700 7514 7512 7404 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01699 7404 7500 7405 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01698 5341 5520 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01697 5429 5813 5341 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01696 4994 5211 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01695 7514 5818 4994 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01694 4994 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01693 7514 5815 4994 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01692 5241 4994 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01691 1468 1419 1338 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01690 1338 1336 1468 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01689 7514 1337 1338 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01688 7514 1310 1308 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01687 1307 1308 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01686 7514 1308 1307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01685 7514 1308 1307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01684 1307 1308 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01683 7514 1310 1311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01682 1309 1311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01681 7514 1311 1309 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01680 7514 1311 1309 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01679 1309 1311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01678 7514 3246 2170 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01677 2169 2170 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01676 7514 2170 2169 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01675 7514 2170 2169 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01674 2169 2170 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01673 7514 3246 2247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01672 2246 2247 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01671 7514 2247 2246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01670 7514 2247 2246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01669 2246 2247 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01668 7514 3246 2248 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01667 2672 2248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01666 7514 2248 2672 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01665 7514 2248 2672 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01664 2672 2248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01663 7514 3246 2178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01662 2177 2178 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01661 7514 2178 2177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01660 7514 2178 2177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01659 2177 2178 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01658 7514 3246 2253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01657 2252 2253 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01656 7514 2253 2252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01655 7514 2253 2252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01654 2252 2253 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01653 7514 3246 2254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01652 2533 2254 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01651 7514 2254 2533 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01650 7514 2254 2533 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01649 2533 2254 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01648 6970 7491 6923 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01647 6923 7379 6970 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01646 7514 7481 6923 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01645 6969 6970 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01644 918 2111 885 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01643 7514 2602 919 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01642 885 919 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01641 2724 3911 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01640 2723 2860 2724 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01639 7514 7420 6072 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01638 6072 6323 6126 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01637 7514 6323 6110 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01636 6126 6110 6073 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01635 6107 6126 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01634 6073 6406 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01633 944 1430 943 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01632 945 1550 944 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01631 943 1688 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01630 1336 944 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01629 7514 1552 945 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01628 945 1867 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01627 7514 3246 3164 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01626 3163 3164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01625 7514 3164 3163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01624 7514 3164 3163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01623 3163 3164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01622 7514 3246 3236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01621 3235 3236 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01620 7514 3236 3235 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01619 7514 3236 3235 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01618 3235 3236 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01617 7514 3246 3237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01616 3581 3237 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01615 7514 3237 3581 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01614 7514 3237 3581 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01613 3581 3237 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01612 7514 3246 3169 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01611 3168 3169 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01610 7514 3169 3168 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01609 7514 3169 3168 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01608 3168 3169 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01607 7514 3246 3245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01606 3244 3245 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01605 7514 3245 3244 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01604 7514 3245 3244 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01603 3244 3245 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01602 7514 3246 3247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01601 3595 3247 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01600 7514 3247 3595 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01599 7514 3247 3595 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01598 3595 3247 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01597 7514 3264 2188 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01596 2187 2188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01595 7514 2188 2187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01594 7514 2188 2187 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01593 2187 2188 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01592 3306 3411 3305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01591 3305 3304 3307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01590 7514 3412 3306 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01589 3303 3307 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01588 4432 6534 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01587 4929 4815 4432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01586 7514 4431 4929 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01585 7514 437 288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01584 602 288 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01583 7514 288 602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01582 7514 288 602 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01581 602 288 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01580 7514 602 395 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01579 5001 395 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01578 7514 395 5001 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01577 7514 395 5001 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01576 5001 395 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01575 7514 602 603 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01574 6133 603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01573 7514 603 6133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01572 7514 603 6133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01571 6133 603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01570 7514 3264 2259 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01569 2260 2259 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01568 7514 2259 2260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01567 7514 2259 2260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01566 2260 2259 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01565 7514 3264 2262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01564 2261 2262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01563 7514 2262 2261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01562 7514 2262 2261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01561 2261 2262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01560 7514 3264 2193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01559 2192 2193 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01558 7514 2193 2192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01557 7514 2193 2192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01556 2192 2193 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01555 7514 3264 2266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01554 2265 2266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01553 7514 2266 2265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01552 7514 2266 2265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01551 2265 2266 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01550 7514 3264 2267 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01549 2553 2267 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01548 7514 2267 2553 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01547 7514 2267 2553 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01546 2553 2267 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01545 7514 3264 3177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01544 3176 3177 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01543 7514 3177 3176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01542 7514 3177 3176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01541 3176 3177 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01540 7514 3264 3254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01539 3253 3254 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01538 7514 3254 3253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01537 7514 3254 3253 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01536 3253 3254 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01535 7514 3264 3255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01534 3466 3255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01533 7514 3255 3466 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01532 7514 3255 3466 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01531 3466 3255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01530 7514 1851 738 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01529 738 2222 763 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01528 762 763 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01527 7514 2157 1928 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01526 1928 1965 1966 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01525 2091 1966 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01524 3513 3922 3512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01523 3512 3925 3513 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01522 7514 5138 3512 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01521 5907 6336 5908 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01520 5908 5905 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01519 5906 6477 5907 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01518 5904 5903 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01517 5903 5902 5906 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01516 7514 5001 3860 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01515 3860 5691 3926 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01514 3925 3926 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01513 6758 6980 6760 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01512 6760 6979 6759 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01511 7514 7464 6758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01510 6757 6759 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01509 4138 4139 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01508 4133 4141 4134 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01507 7514 4933 4133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01506 7514 4277 4141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01505 4140 4141 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01504 7514 4572 4139 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01503 4135 4136 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01502 7514 4135 4137 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01501 4134 4140 4135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01500 4933 4134 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01499 7514 4134 4933 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01498 4137 4140 4136 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01497 4136 4141 4138 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01496 6732 6965 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01495 4361 4933 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01494 2589 3418 2588 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01493 2588 2929 2589 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01492 7514 6035 2588 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01491 3841 5001 3842 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01490 3842 5691 3843 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01489 7514 5690 3841 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01488 3840 3843 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01487 6899 7227 6900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01486 6900 7228 6899 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01485 7514 7475 6900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01484 3724 3890 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01483 7173 7387 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01482 7369 7480 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01481 6671 7045 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01480 6713 6991 6671 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01479 7514 5092 4825 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01478 4825 5716 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01477 7514 4824 4825 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01476 6595 6682 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01475 6594 6593 6595 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01474 1204 2255 1205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01473 1205 1369 1204 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01472 7514 4161 1205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01471 1570 1204 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01470 1510 1631 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01469 1979 1581 1510 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01468 7514 3184 3185 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01467 3185 3356 3186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01466 3183 3186 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01465 6452 7033 6454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01464 6453 7267 6452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01463 6454 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01462 6451 6452 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01461 7514 7032 6453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01460 6453 7137 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01459 1614 1898 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01458 1753 1688 1614 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01457 5169 5523 5168 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01456 5168 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01455 5167 5841 5169 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01454 5166 5690 5167 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01453 6608 6342 6343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01452 6343 6340 6608 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01451 7514 6341 6343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01450 5091 5378 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01449 7514 6910 5091 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01448 5091 6981 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01447 7514 5377 5091 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01446 5087 5091 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01445 7514 5882 4417 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01444 4417 4912 4419 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01443 7514 4912 4420 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01442 4419 4420 4418 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01441 4416 4419 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01440 4418 5138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01439 7514 6025 4177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01438 4177 4912 4202 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01437 7514 4912 4203 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01436 4202 4203 4178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01435 4475 4202 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01434 4178 5137 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01433 4851 5071 4850 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01432 4850 4847 4849 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01431 7514 4848 4851 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01430 4846 4849 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01429 3044 3081 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01428 3082 3226 3044 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01427 7514 324 325 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01426 324 1851 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01425 325 2708 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01424 2172 4568 2173 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01423 2173 2185 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01422 3214 2171 2172 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01421 7514 4983 4982 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01420 4983 5291 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01419 4982 5365 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01418 4764 6030 4613 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01417 4613 6029 4764 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01416 7514 5069 4613 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01415 5480 7018 5479 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01414 5479 5521 5522 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01413 7514 5816 5480 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01412 5520 5522 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01411 2642 2687 2641 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01410 2641 2684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01409 2685 4000 2642 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01408 7514 2655 2651 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01407 7514 2648 2651 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01406 2651 2647 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01405 6165 2651 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01404 5938 6112 5939 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01403 5939 6336 5993 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01402 7514 6576 5938 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01401 5992 5993 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01400 1417 1813 1391 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01399 1390 1679 1417 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01398 1391 1684 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01397 1473 1417 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01396 7514 1680 1390 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01395 1390 1681 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01394 7514 908 743 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01393 743 828 774 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01392 1032 774 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01391 7514 2522 2524 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01390 2522 2521 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01389 2524 3239 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01388 6957 7496 6928 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01387 6928 7289 6957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01386 7514 6981 6928 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01385 3145 3214 3146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01384 3146 3212 3145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01383 7514 3879 3146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01382 7514 5889 4146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01381 4146 4724 4147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01380 4224 4147 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01379 2995 2543 2036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01378 2036 2541 2995 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01377 7514 2035 2036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01376 452 500 685 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01375 7514 939 452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01374 453 762 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01373 685 499 453 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01372 7514 762 500 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01371 499 939 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01370 733 4442 732 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01369 732 1051 734 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01368 7514 2880 733 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01367 731 734 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01366 7514 4376 4162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01365 4162 4161 4163 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01364 5172 4163 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01363 7514 4600 1245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01362 1245 2033 1313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01361 1312 1313 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01360 3849 3886 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01359 3847 3888 3881 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01358 7514 3879 3847 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01357 7514 4488 3888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01356 3889 3888 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01355 7514 3884 3886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01354 3883 3885 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01353 7514 3883 3848 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01352 3881 3889 3883 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01351 3879 3881 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01350 7514 3881 3879 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01349 3848 3889 3885 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01348 3885 3888 3849 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01347 4981 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01346 5364 7286 4981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01345 4980 4979 5364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01344 7514 5275 4980 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01343 4980 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01342 15 16 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01341 10 18 11 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01340 7514 5125 10 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01339 7514 360 18 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01338 17 18 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01337 7514 5124 16 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01336 12 13 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01335 7514 12 14 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01334 11 17 12 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01333 5125 11 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01332 7514 11 5125 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01331 14 17 13 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01330 13 18 15 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01329 7514 4411 4414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01328 4414 4412 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01327 4410 4415 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01326 4414 4413 4415 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01325 4415 4916 4414 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_01324 4191 4447 4192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01323 4192 4448 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01322 4190 4442 4191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01321 5842 4235 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01320 4235 4934 4190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01319 7039 7227 7040 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01318 7040 7228 7039 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01317 7514 7480 7040 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01316 7514 6653 6912 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01315 6653 7384 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01314 6912 6852 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01313 7514 4995 4932 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01312 4932 4996 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01311 5273 4932 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01310 2987 4359 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01309 2986 3097 2987 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01308 7514 6944 5028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01307 5028 5072 5073 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01306 5071 5073 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01305 227 518 226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01304 226 283 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01303 514 225 227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01302 617 640 616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01301 616 1029 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01300 615 1145 617 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01299 641 1809 615 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01298 7264 7309 7265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01297 7265 7416 7264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01296 7514 7420 7265 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01295 7514 7354 6508 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01294 6508 6576 6575 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01293 6535 6575 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01292 4817 6534 4818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01291 4818 5226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01290 4816 4829 4817 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01289 5072 4864 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01288 4864 4815 4816 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01287 2342 2418 2368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01286 2368 2789 2343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01285 2343 2505 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01284 2341 2504 2368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01283 7514 2416 2341 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01282 7514 2502 2342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01281 2366 2368 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01280 7514 1688 349 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01279 349 1082 379 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01278 378 379 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01277 1944 1976 1945 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01276 1945 2591 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01275 1943 3820 1944 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01274 2542 1977 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01273 1977 4376 1943 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01272 1805 4600 1804 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01271 1804 4603 1839 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01270 7514 7042 1805 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01269 1838 1839 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01268 4546 4547 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01267 4542 4548 4541 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01266 7514 4975 4542 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01265 7514 4638 4548 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01264 4549 4548 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01263 7514 4641 4547 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01262 4543 4545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01261 7514 4543 4544 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01260 4541 4549 4543 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01259 4975 4541 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01258 7514 4541 4975 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01257 4544 4549 4545 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01256 4545 4548 4546 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01255 4290 4448 4291 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01254 4291 4441 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01253 4288 5173 4290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01252 5718 4289 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01251 4289 4446 4288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01250 1251 1384 1252 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01249 1252 2392 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01248 1250 3820 1251 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01247 1574 1298 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01246 1298 2881 1250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01245 4143 4069 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01244 7196 7453 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01243 7455 7454 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01242 5082 5376 4993 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01241 4993 5273 5082 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01240 7514 6035 4993 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01239 7514 4579 4274 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01238 7514 4774 4274 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01237 4274 5069 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01236 4715 4274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01235 5366 5735 5340 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01234 5340 5734 5366 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01233 7514 5815 5340 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01232 6323 7494 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01231 6770 7108 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01230 2753 2889 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01229 2752 2751 2753 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01228 166 446 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01227 233 3248 166 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01226 133 239 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01225 132 4296 133 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01224 7514 6386 6307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01223 6307 6306 6308 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01222 6310 6308 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01221 6210 6632 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01220 6825 6242 6210 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01219 4910 4908 4876 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01218 4876 5369 4910 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01217 7514 5226 4876 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01216 5660 4910 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01215 7514 6386 6353 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01214 6353 6389 6387 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01213 6633 6387 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01212 7514 6175 4706 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01211 4706 4912 4707 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01210 7514 4912 4708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01209 4707 4708 4709 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01208 4705 4707 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01207 4709 4834 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01206 7514 5887 3785 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01205 3785 4912 3787 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01204 7514 4912 3788 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01203 3787 3788 3786 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01202 4040 3787 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01201 3786 5274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01200 251 1082 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01199 275 1688 251 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01198 3139 3403 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01197 3138 3137 3139 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01196 347 2696 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01195 509 1851 347 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01194 2364 5841 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01193 2395 5840 2364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01192 2363 2398 2395 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01191 7514 2540 2363 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01190 2362 2536 2395 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01189 7514 2684 2362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01188 3633 3069 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01187 7514 3070 3633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01186 3633 3071 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01185 7514 3074 3633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01184 5490 5539 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01183 5540 5667 5490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01182 5717 5904 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01181 5716 5891 5717 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01180 3062 3119 3063 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01179 3063 3351 3118 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01178 7514 3266 3062 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01177 3181 3118 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01176 7514 6035 4711 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01175 4711 4912 4712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01174 7514 4912 4714 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01173 4712 4714 4713 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01172 4710 4712 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01171 4713 5043 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01170 2662 2945 2440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01169 2440 2946 2662 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01168 7514 5216 2440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01167 5786 7042 5785 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01166 5785 6332 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01165 5844 7162 5786 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01164 7514 1037 650 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01163 650 2300 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01162 775 650 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01161 2659 2229 2058 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01160 2058 2154 2659 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01159 7514 2164 2058 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01158 4584 4582 4586 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01157 4586 4585 4587 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01156 7514 4583 4584 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01155 4581 4587 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01154 7514 6846 6769 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01153 6769 6770 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01152 6768 6769 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01151 346 365 6168 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01150 7514 363 346 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01149 345 558 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01148 6168 362 345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01147 7514 558 365 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01146 362 363 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01145 4886 4933 4887 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01144 4887 5718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01143 4885 5001 4886 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01142 6131 4934 4885 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01141 1248 1809 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01140 2027 1954 1248 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01139 1247 1339 2027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01138 7514 1266 1247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01137 1247 1267 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_01136 1393 1813 1392 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01135 1392 1420 1421 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01134 7514 1556 1393 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01133 1419 1421 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01132 6712 6770 6670 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01131 6670 6846 6712 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01130 7514 7354 6670 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01129 6710 6712 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01128 4457 4489 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01127 4455 4491 4484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01126 7514 6035 4455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01125 7514 4488 4491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01124 4490 4491 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01123 7514 4710 4489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01122 4483 4486 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01121 7514 4483 4456 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01120 4484 4490 4483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01119 6035 4484 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01118 7514 4484 6035 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01117 4456 4490 4486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01116 4486 4491 4457 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01115 3374 3820 3966 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01114 7514 3820 3422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01113 3375 3819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01112 3966 3422 3375 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01111 7514 3993 3374 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01110 7514 5686 6394 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01109 5686 6333 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01108 6394 5685 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01107 4311 4344 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01106 4309 4346 4339 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01105 7514 6175 4309 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01104 7514 4638 4346 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01103 4345 4346 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_01102 7514 4705 4344 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_01101 4341 4342 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01100 7514 4341 4310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01099 4339 4345 4341 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01098 6175 4339 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01097 7514 4339 6175 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01096 4310 4345 4342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01095 4342 4346 4311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01094 1890 2171 1889 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01093 1889 2318 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01092 1888 2102 1890 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01091 4413 1887 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01090 1887 4773 1888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01089 1673 4377 1674 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01088 1674 1707 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01087 1672 5173 1673 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01086 1833 1708 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_01085 1708 4376 1672 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01084 7514 1023 936 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01083 936 1022 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01082 7514 1021 936 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01081 6207 6236 6234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01080 7514 6629 6207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01079 6208 6553 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01078 6234 6233 6208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01077 7514 6553 6236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01076 6233 6629 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01075 3741 3739 3689 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01074 3689 3738 3741 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01073 7514 3736 3689 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01072 3737 3741 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01071 4308 5826 4307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01070 4307 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01069 4701 6539 4308 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01068 7365 7362 7366 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01067 7514 7475 7365 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01066 7364 7471 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01065 7366 7363 7364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01064 7514 7471 7362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01063 7363 7475 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01062 7514 2109 2183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01061 2183 2042 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01060 7514 2328 2183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01059 2870 3179 2871 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01058 2871 2869 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01057 2868 2954 2870 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01056 3109 2995 2868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01055 6356 6968 6355 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01054 6355 6967 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01053 6391 7494 6356 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01052 50 82 225 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01051 7514 186 50 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01050 51 325 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01049 225 81 51 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01048 7514 325 82 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01047 81 186 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01046 4442 1449 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01045 7514 1168 4442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01044 4442 2111 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01043 7514 2602 4442 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01042 3369 4367 3370 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01041 3370 4368 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01040 3368 4985 3369 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01039 3418 6408 3368 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01038 1142 1430 1117 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01037 1116 1332 1142 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01036 1117 3546 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01035 1464 1142 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01034 7514 1333 1116 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01033 1116 1334 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_01032 6554 7491 6499 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01031 6499 7379 6554 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01030 7514 6676 6499 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01029 6523 6554 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01028 5607 5606 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01027 7514 5818 5607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01026 5607 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01025 7514 5815 5607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_01024 5828 5607 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01023 7514 4296 4298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01022 4298 5251 4299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01021 4297 4299 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01020 1118 1144 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01019 1258 1342 1118 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01018 6681 5735 5736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01017 5736 5734 6681 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01016 7514 6315 5736 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01015 4926 5376 4881 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01014 4881 5273 4926 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01013 7514 6175 4881 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_01012 7514 3993 3818 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01011 3818 3820 3822 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01010 7514 3820 3823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01009 3822 3823 3821 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01008 3817 3822 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01007 3821 3819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_01006 3175 4600 3174 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01005 3174 4603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01004 3173 6133 3175 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01003 4724 6333 3173 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_01002 6727 7452 6728 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01001 6728 7074 6729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_01000 7514 7453 6727 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00999 6726 6729 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00998 1122 1341 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00997 7514 1342 1122 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00996 1122 1270 1153 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00995 1153 1866 1122 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00994 7514 6846 5622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00993 5622 5619 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00992 5685 5621 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00991 5622 5620 5621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00990 5621 6770 5622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00989 7514 2836 2623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00988 2623 2841 2646 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00987 2645 2646 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00986 1901 2816 1900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00985 1900 2454 1901 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00984 7514 1899 1900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00983 1898 1901 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00982 7514 2657 2625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00981 2625 3213 2656 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00980 2705 2656 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00979 3026 3029 3028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00978 3028 3033 3027 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00977 7514 3030 3026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00976 3663 3027 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00975 7514 5171 4189 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00974 4189 5172 4234 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00973 4603 4234 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00972 1637 1676 3412 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00971 7514 1858 1637 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00970 1638 1954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00969 3412 1677 1638 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00968 7514 1954 1676 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00967 1677 1858 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00966 3852 3897 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00965 3850 3900 3893 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00964 7514 3890 3850 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00963 7514 4561 3900 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00962 3899 3900 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00961 7514 3895 3897 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00960 3894 3896 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00959 7514 3894 3851 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00958 3893 3899 3894 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00957 3890 3893 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00956 7514 3893 3890 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00955 3851 3899 3896 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00954 3896 3900 3852 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00953 6845 5001 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00952 3427 4148 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00951 7514 4996 4823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00950 4823 4822 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00949 7514 7227 4823 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00948 3537 3593 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00947 3535 3596 3586 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00946 7514 3997 3535 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00945 7514 3595 3596 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00944 3594 3596 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00943 7514 3592 3593 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00942 3588 3590 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00941 7514 3588 3536 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00940 3586 3594 3588 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00939 3997 3586 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00938 7514 3586 3997 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00937 3536 3594 3590 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00936 3590 3596 3537 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00935 3665 4156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00934 1709 1906 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00933 4593 5841 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00932 1134 1620 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00931 1572 1619 1134 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00930 980 1575 981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00929 981 978 980 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00928 7514 1106 981 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00927 979 980 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00926 4071 4282 4022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00925 4022 4360 4071 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00924 7514 6703 4022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00923 4070 4071 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00922 7103 7334 7038 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00921 7038 7383 7103 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00920 7514 7452 7038 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00919 6597 6598 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00918 6750 6596 6597 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00917 3136 3135 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00916 3134 3644 3136 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00915 1641 1732 1516 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00914 1516 1547 1641 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00913 7514 1548 1516 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00912 4400 4673 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00911 7283 4674 4400 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00910 7514 4756 4758 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00909 4756 4755 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00908 4758 4754 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00907 5156 5376 5033 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00906 5033 5273 5156 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00905 7514 6392 5033 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00904 6322 6323 6321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00903 6321 6406 6322 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00902 7514 7420 6321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00901 7514 3820 867 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00900 867 6344 914 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00899 7514 6344 888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00898 914 888 868 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00897 915 914 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00896 868 5138 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00895 7514 4158 590 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00894 590 6344 658 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00893 7514 6344 660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00892 658 660 591 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00891 656 658 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00890 591 5137 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00889 7514 1168 842 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00888 842 6344 869 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00887 7514 6344 870 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00886 869 870 843 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00885 841 869 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00884 843 5216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00883 1194 1968 1195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00882 1195 2718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00881 1193 1700 1194 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00880 1341 1688 1193 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00879 3688 3732 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00878 5616 3733 3688 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00877 3687 3734 5616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00876 7514 3967 3687 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00875 3686 3920 5616 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00874 7514 4077 3686 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00873 4601 4603 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00872 4602 4600 4601 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00871 1148 1146 1119 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00870 1119 1182 1148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00869 7514 1145 1119 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00868 1954 1148 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00867 4591 4588 4590 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00866 4590 4667 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00865 4821 4589 4591 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00864 7514 2602 2604 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00863 2604 6344 2606 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00862 7514 6344 2607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00861 2606 2607 2605 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00860 2603 2606 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00859 2605 5055 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00858 7514 483 1775 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00857 483 4376 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00856 1775 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00855 1372 2543 1237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00854 1237 2541 1372 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00853 7514 1628 1237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00852 1894 1893 1895 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00851 1895 2104 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00850 1891 1896 1894 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00849 1892 6407 1891 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00848 5451 6565 5452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00847 5452 6566 5451 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00846 7514 7454 5452 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00845 983 2392 984 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00844 984 1976 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00843 982 3820 983 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00842 1441 4376 982 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00841 5811 5885 5598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00840 5598 5884 5811 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00839 7514 6125 5598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00838 1626 1709 1625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00837 1625 1624 1626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00836 7514 4597 1625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00835 1899 1626 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00834 6247 6393 5888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00833 5888 6394 6247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00832 7514 5887 5888 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00831 7514 3352 1200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00830 1200 1577 1229 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00829 2504 1229 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00828 4272 4367 4271 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00827 4271 4368 4273 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00826 7514 4985 4272 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00825 4566 4273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00824 6086 6708 6085 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00823 6085 6131 6130 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00822 7514 6533 6086 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00821 6705 6130 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00820 3679 4588 3680 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00819 3680 4568 3716 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00818 7514 4569 3679 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00817 4411 3716 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00816 3862 4069 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00815 7432 4228 3862 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00814 3861 4378 7432 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00813 7514 4149 3861 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00812 3861 5909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00811 5460 6652 5321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00810 5321 5467 5460 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00809 7514 7235 5321 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00808 3048 3094 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00807 3046 3096 3088 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00806 7514 3086 3046 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00805 7514 3571 3096 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00804 3095 3096 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00803 7514 3092 3094 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00802 3089 3091 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00801 7514 3089 3047 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00800 3088 3095 3089 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00799 3086 3088 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00798 7514 3088 3086 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00797 3047 3095 3091 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00796 3091 3096 3048 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00795 6976 6894 6895 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00794 6895 6893 6976 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00793 7514 6892 6895 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00792 4195 6168 4176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00791 4176 6169 4195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00790 7514 5069 4176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00789 274 3081 250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00788 250 2134 274 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00787 7514 272 250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00786 699 274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00785 7298 7332 7317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00784 7514 7494 7298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00783 7299 7493 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00782 7317 7333 7299 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00781 7514 7493 7332 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00780 7333 7494 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00779 6482 6489 6483 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00778 6481 6490 6482 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00777 6491 6482 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00776 7514 6482 6491 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00775 6487 6488 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00774 7514 6613 6488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00773 6489 6490 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00772 7514 6611 6490 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00771 6484 6486 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00770 6483 7500 6484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00769 6486 6490 6487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00768 6485 6489 6486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00767 7514 6483 6485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00766 7514 6491 6480 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00765 6480 7500 6481 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00764 3292 3293 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00763 3288 3295 3287 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00762 7514 3475 3288 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00761 7514 3400 3295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00760 3294 3295 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00759 7514 3476 3293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00758 3289 3290 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00757 7514 3289 3291 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00756 3287 3294 3289 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00755 3475 3287 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00754 7514 3287 3475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00753 3291 3294 3290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00752 3290 3295 3292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00751 2620 2543 1950 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00750 1950 2541 2620 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00749 7514 1979 1950 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00748 4832 5826 4831 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00747 4831 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00746 4833 5045 4832 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00745 6966 7033 6935 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00744 6934 7016 6966 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00743 6935 7034 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00742 6944 6966 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00741 7514 7032 6934 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00740 6934 7307 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00739 826 3546 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00738 827 1430 826 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00737 825 900 827 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00736 7514 823 825 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00735 825 824 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00734 431 3546 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00733 467 2016 431 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00732 7514 647 467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00731 464 467 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00730 1070 2139 1069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00729 1069 3545 1070 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00728 7514 1688 1069 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00727 1068 1070 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00726 3660 4084 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00725 7514 4006 3660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00724 3660 3840 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00723 7514 3927 3660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00722 5484 5677 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00721 5535 5534 5484 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00720 2352 2862 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00719 2435 2589 2352 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00718 7514 1699 1485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00717 1485 3159 1486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00716 7514 3159 1487 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00715 1486 1487 1488 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00714 1746 1486 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00713 1488 1883 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.67U AS=0.1742P AD=0.1742P PS=1.87U PD=1.87U 
Mtr_00712 2782 3119 2783 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00711 2783 2825 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00710 2781 3266 2782 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00709 2971 3814 2781 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00708 4836 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00707 4837 7286 4836 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00706 4835 4834 4837 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00705 7514 5275 4835 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00704 4835 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00703 6044 7227 6045 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00702 6045 7228 6044 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00701 7514 7494 6045 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00700 3548 3549 3519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00699 3519 3545 3548 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00698 7514 3546 3519 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00697 7514 7480 7397 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00696 7397 7477 7423 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00695 7471 7423 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00694 5002 5001 5003 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00693 5003 5718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00692 6708 5000 5002 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00691 363 893 315 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00690 315 455 363 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00689 7514 641 315 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00688 707 706 708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00687 708 709 707 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00686 7514 1342 708 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00685 6030 707 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00684 4434 6133 4435 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00683 4435 4728 4436 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00682 7514 6333 4434 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00681 4996 4436 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00680 5731 5728 5730 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00679 5730 6378 5732 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00678 7514 5729 5731 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00677 5727 5732 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00676 5023 7164 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00675 5056 7286 5023 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00674 5022 5055 5056 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00673 7514 5275 5022 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00672 5022 5273 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00671 7514 5451 5164 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00670 5164 5166 5165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00669 5306 5165 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00668 7514 2685 2464 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00667 2464 2465 2466 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00666 2463 2466 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00665 7400 7489 7399 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00664 7399 7481 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00663 7398 7493 7400 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00662 7477 7425 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00661 7425 7494 7398 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00660 60 108 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00659 58 110 102 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00658 7514 1906 58 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00657 7514 403 110 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00656 109 110 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00655 7514 132 108 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00654 104 105 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00653 7514 104 59 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00652 102 109 104 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00651 1906 102 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00650 7514 102 1906 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00649 59 109 105 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00648 105 110 60 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00647 4921 5376 4737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00646 4737 5273 4921 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00645 7514 6025 4737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00644 7514 1466 1083 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00643 1083 1430 1084 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00642 3545 1084 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00641 7514 3483 3486 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00640 3486 3484 3485 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00639 3482 3485 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00638 7514 1767 1769 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00637 1769 2395 1770 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00636 1768 1770 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00635 1568 2255 1364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00634 1364 1363 1568 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00633 7514 1449 1364 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00632 7514 1111 756 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00631 756 1112 795 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00630 1047 795 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00629 7065 7103 7066 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00628 7066 7105 7106 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00627 7514 7156 7065 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00626 7104 7106 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00625 6084 6980 6083 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00624 6083 6979 6127 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00623 7514 7466 6084 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00622 6111 6127 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00621 729 918 445 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00620 445 481 729 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00619 7514 3427 445 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00618 3684 3727 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00617 5835 4228 3684 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00616 3683 3819 5835 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00615 7514 4149 3683 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00614 3683 5909 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00613 243 4437 245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00612 245 4081 244 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00611 7514 5001 243 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00610 242 244 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00609 205 208 1633 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00608 7514 890 205 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00607 207 1736 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00606 1633 206 207 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00605 7514 1736 208 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00604 206 890 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00603 5146 5147 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00602 5142 5149 5141 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00601 7514 5833 5142 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00600 7514 5518 5149 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00599 5148 5149 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00598 7514 5229 5147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00597 5143 5144 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00596 7514 5143 5145 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00595 5141 5148 5143 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00594 5833 5141 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00593 7514 5141 5833 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00592 5145 5148 5144 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00591 5144 5149 5146 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00590 2255 2602 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00589 2103 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00588 5000 4934 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00587 171 1021 165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00586 165 1022 171 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00585 7514 1023 165 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00584 937 171 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00583 1395 1435 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00582 1422 1768 1395 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00581 1394 1556 1422 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00580 7514 1682 1394 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00579 1394 1479 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.95U AS=0.507P AD=0.507P PS=4.42U PD=4.42U 
Mtr_00578 1509 1508 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00577 4296 7162 1509 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00576 6626 6623 6625 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00575 7514 6732 6626 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00574 6627 6869 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00573 6625 6624 6627 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00572 7514 6869 6623 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00571 6624 6732 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00570 6465 6697 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00569 6466 6464 6465 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00568 5329 7390 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00567 6135 6652 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00566 4751 4780 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00565 4822 4781 4751 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00564 6034 6032 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00563 6690 6033 6034 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00562 5668 5653 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00561 7514 5818 5668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00560 5668 5819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00559 7514 5815 5668 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00558 5669 5668 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00557 830 828 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00556 829 908 830 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00555 7068 7109 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00554 7110 7108 7068 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00553 3042 3482 3043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00552 3043 3080 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00551 3143 3079 3042 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00550 1402 1883 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00549 1567 1699 1402 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00548 4467 4569 4466 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00547 4466 4568 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00546 4820 4773 4467 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00545 2032 4600 2034 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00544 2034 2033 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00543 4726 7162 2032 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00542 2199 2524 2198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00541 2198 4694 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00540 2418 2228 2199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00539 6033 6030 6031 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00538 6031 6029 6033 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00537 7514 6315 6031 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00536 4019 4368 4020 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00535 4020 5085 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00534 4018 4367 4019 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00533 5069 4985 4018 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00532 2256 2543 2043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00531 2043 2541 2256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00530 7514 2179 2043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00529 2921 2958 2920 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00528 2920 2988 2957 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00527 7514 2956 2921 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00526 6046 2957 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00525 5154 5274 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00524 5300 5832 5154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00523 7514 5153 5300 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00522 2657 3418 2348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00521 2348 2929 2657 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00520 7514 6392 2348 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00519 7514 4082 4447 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00518 4082 4158 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00517 4447 4161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00516 6059 6114 6060 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00515 6060 6535 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00514 6057 6773 6059 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00513 6058 6056 6057 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00512 4620 4659 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00511 4618 4662 4654 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00510 7514 5454 4618 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00509 7514 4660 4662 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00508 4661 4662 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00507 7514 4779 4659 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00506 4655 4658 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00505 7514 4655 4619 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00504 4654 4661 4655 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00503 5454 4654 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00502 7514 4654 5454 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00501 4619 4661 4658 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00500 4658 4662 4620 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00499 2136 2286 2135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00498 2135 3131 2136 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00497 7514 2133 2135 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00496 2134 2136 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00495 3469 936 938 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00494 938 937 3469 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00493 7514 1342 938 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00492 3719 3501 3008 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00491 3008 4669 3719 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00490 7514 3226 3008 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00489 3645 4431 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00488 3226 4991 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00487 890 2095 850 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00486 850 3545 890 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00485 7514 1688 850 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00484 3917 3545 1094 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00483 1094 2027 3917 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00482 7514 2029 1094 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00481 3646 4718 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00480 3012 4424 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00479 4378 4937 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00478 754 1441 755 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00477 755 1236 794 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00476 7514 844 754 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00475 978 794 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00474 7514 1775 482 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00473 482 1052 537 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00472 536 537 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00471 5581 6894 5475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00470 5475 5902 5581 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00469 7514 5507 5475 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00468 586 588 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00467 581 589 580 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00466 7514 579 581 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00465 7514 788 589 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00464 587 589 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00463 7514 584 588 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00462 582 585 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00461 7514 582 583 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00460 580 587 582 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00459 579 580 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00458 7514 580 579 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00457 583 587 585 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00456 585 589 586 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00455 3404 3481 3362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00454 3362 4695 3404 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00453 7514 3484 3362 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00452 3403 3404 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00451 1071 1952 1073 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00450 1072 1337 1071 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00449 1073 1548 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00448 1074 1071 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00447 7514 1419 1072 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00446 1072 1336 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00445 4009 4043 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00444 4007 4044 4037 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00443 7514 5887 4007 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00442 7514 4638 4044 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00441 4045 4044 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00440 7514 4040 4043 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00439 4039 4042 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00438 7514 4039 4008 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00437 4037 4045 4039 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00436 5887 4037 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00435 7514 4037 5887 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00434 4008 4045 4042 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00433 4042 4044 4009 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00432 290 297 292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00431 258 298 290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00430 4376 290 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00429 7514 290 4376 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00428 261 296 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00427 7514 295 296 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00426 297 298 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00425 7514 403 298 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00424 260 294 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00423 292 7500 260 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00422 294 298 261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00421 259 297 294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00420 7514 292 259 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00419 7514 4376 257 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00418 257 7500 258 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00417 6318 6393 6176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00416 6176 6394 6318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00415 7514 6175 6176 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00414 405 242 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00413 7514 195 405 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00412 7514 4821 4777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00411 4777 4819 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00410 7514 4820 4777 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00409 2763 2854 2802 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00408 2802 2800 2764 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00407 2764 2801 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00406 2762 2991 2802 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00405 7514 2995 2762 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00404 7514 4410 2763 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00403 2798 2802 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00402 3918 5889 3859 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00401 3859 3917 3918 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00400 7514 4825 3859 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00399 4075 3918 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00398 5333 5826 5332 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00397 5332 5351 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00396 5498 5350 5333 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00395 941 2222 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00394 942 1851 941 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00393 1554 1552 1517 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00392 1517 1867 1554 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00391 7514 1550 1517 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00390 1551 1554 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00389 6877 6878 6880 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00388 6880 7264 6879 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00387 7514 6947 6877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00386 6876 6879 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00385 7514 5299 5301 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00384 5301 5300 5302 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00383 5438 5302 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00382 2792 3481 2759 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00381 2759 4695 2792 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00380 7514 3077 2759 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00379 6763 7104 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00378 6762 6761 6763 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00377 7514 5312 4223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00376 4222 4223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00375 7514 4223 4222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00374 7514 4223 4222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00373 4222 4223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00372 7514 5312 4276 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00371 4275 4276 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00370 7514 4276 4275 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00369 7514 4276 4275 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00368 4275 4276 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00367 7514 5312 4278 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00366 4277 4278 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00365 7514 4278 4277 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00364 7514 4278 4277 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00363 4277 4278 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00362 7514 5312 4227 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00361 4226 4227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00360 7514 4227 4226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00359 7514 4227 4226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00358 4226 4227 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00357 7514 5312 4284 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00356 4283 4284 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00355 7514 4284 4283 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00354 7514 4284 4283 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00353 4283 4284 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00352 7514 5312 4285 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00351 4660 4285 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00350 7514 4285 4660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00349 7514 4285 4660 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00348 4660 4285 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00347 7514 5312 5240 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00346 5239 5240 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00345 7514 5240 5239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00344 7514 5240 5239 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00343 5239 5240 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00342 314 1680 313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00341 313 1681 314 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00340 7514 1679 313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00339 312 314 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00338 1780 1810 1781 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00337 1781 1954 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00336 2008 1809 1780 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00335 2621 2620 2622 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00334 2622 4524 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00333 2619 3431 2621 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00332 2618 2823 2619 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00331 7514 269 455 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00330 269 462 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00329 455 1021 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00328 2994 3137 2992 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00327 2992 2991 2993 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00326 2993 2995 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00325 2990 3082 2992 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00324 7514 3701 2990 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00323 7514 3403 2994 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00322 3406 2992 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00321 1345 1340 1344 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00320 1343 1341 1345 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00319 1344 1342 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00318 1339 1345 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00317 7514 1551 1343 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00316 1343 1741 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00315 7514 5312 5304 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00314 5303 5304 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00313 7514 5304 5303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00312 7514 5304 5303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00311 5303 5304 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00310 7514 5312 5305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00309 5531 5305 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00308 7514 5305 5531 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00307 7514 5305 5531 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00306 5531 5305 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00305 7514 5312 5246 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00304 5245 5246 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00303 7514 5246 5245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00302 7514 5246 5245 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00301 5245 5246 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00300 7514 5312 5311 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00299 5310 5311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00298 7514 5311 5310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00297 7514 5311 5310 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00296 5310 5311 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00295 7514 5312 5313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00294 5449 5313 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00293 7514 5313 5449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00292 7514 5313 5449 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00291 5449 5313 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00290 7514 5327 4233 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00289 4232 4233 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00288 7514 4233 4232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00287 7514 4233 4232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00286 4232 4233 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00285 7514 5327 4293 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00284 4292 4293 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00283 7514 4293 4292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00282 7514 4293 4292 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00281 4292 4293 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00280 7514 5327 4295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00279 4294 4295 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00278 7514 4295 4294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00277 7514 4295 4294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00276 4294 4295 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00275 7514 1851 1737 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00274 1737 1876 1738 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00273 1736 1738 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00272 2916 3160 2917 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00271 2917 3303 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00270 2915 3159 2916 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00269 2951 2952 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.87U AS=0.4862P AD=0.4862P PS=4.27U PD=4.27U 
Mtr_00268 2952 3326 2915 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00267 6162 6234 6161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00266 6161 6160 6162 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00265 7514 7420 6161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00264 7514 2836 2838 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00263 2838 3128 2839 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00262 2837 2839 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00261 6473 6565 6472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00260 6472 6566 6473 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00259 7514 7335 6472 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00258 7514 5327 4237 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00257 4236 4237 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00256 7514 4237 4236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00255 7514 4237 4236 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00254 4236 4237 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00253 7514 5327 4304 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00252 4303 4304 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00251 7514 4304 4303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00250 7514 4304 4303 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00249 4303 4304 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00248 7514 5327 4306 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00247 4305 4306 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00246 7514 4306 4305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00245 7514 4306 4305 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00244 4305 4306 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00243 7514 5327 5248 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00242 5247 5248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00241 7514 5248 5247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00240 7514 5248 5247 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00239 5247 5248 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00238 7514 5327 5318 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00237 5317 5318 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00236 7514 5318 5317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00235 7514 5318 5317 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00234 5317 5318 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00233 7514 5327 5320 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00232 5319 5320 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00231 7514 5320 5319 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00230 7514 5320 5319 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00229 5319 5320 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00228 7514 5327 5255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00227 5254 5255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00226 7514 5255 5254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00225 7514 5255 5254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00224 5254 5255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00223 7514 2657 2480 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00222 2480 2856 2509 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00221 2846 2509 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00220 341 340 342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00219 342 399 341 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00218 7514 5619 342 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00217 1109 341 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00216 1606 1883 1608 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00215 1607 3546 1606 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00214 1608 1851 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00213 1605 1606 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00212 7514 1823 1607 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00211 1607 3545 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00210 1877 2424 1879 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00209 1879 1876 1878 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00208 7514 2220 1877 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00207 2093 1878 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00206 7290 7324 7307 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00205 7514 7462 7290 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00204 7291 7413 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00203 7307 7325 7291 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00202 7514 7413 7324 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00201 7325 7462 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00200 574 1155 573 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00199 573 775 575 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00198 7514 1688 574 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00197 653 575 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00196 1000 1968 1001 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00195 1001 2718 1036 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00194 7514 1700 1000 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00193 1430 1036 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.17U AS=0.5642P AD=0.5642P PS=4.87U PD=4.87U 
Mtr_00192 2030 5889 2031 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00191 2028 2029 2030 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00190 2031 4568 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00189 2820 2030 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00188 7514 3545 2028 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00187 2028 2027 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.1U AS=0.546P AD=0.546P PS=4.72U PD=4.72U 
Mtr_00186 7514 5327 5326 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00185 5325 5326 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00184 7514 5326 5325 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00183 7514 5326 5325 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00182 5325 5326 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00181 7514 5327 5328 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00180 5554 5328 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00179 7514 5328 5554 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00178 7514 5328 5554 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00177 5554 5328 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00176 7514 7224 6178 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00175 6177 6178 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00174 7514 6178 6177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00173 7514 6178 6177 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00172 6177 6178 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00171 7514 7224 6250 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00170 6249 6250 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00169 7514 6250 6249 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00168 7514 6250 6249 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00167 6249 6250 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00166 7514 7224 6251 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00165 6693 6251 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00164 7514 6251 6693 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00163 7514 6251 6693 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00162 6693 6251 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00161 7514 7224 6184 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00160 6183 6184 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00159 7514 6184 6183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00158 7514 6184 6183 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00157 6183 6184 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00156 7514 7224 6255 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00155 6254 6255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00154 7514 6255 6254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00153 7514 6255 6254 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00152 6254 6255 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00151 7514 7224 6257 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00150 6256 6257 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00149 7514 6257 6256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00148 7514 6257 6256 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00147 6256 6257 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00146 3985 3987 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00145 3959 3988 3984 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00144 7514 4215 3959 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00143 7514 4277 3988 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00142 3986 3988 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.05U AS=0.273P AD=0.273P PS=2.62U PD=2.62U 
Mtr_00141 7514 4216 3987 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.35U AS=0.351P AD=0.351P PS=3.22U PD=3.22U 
Mtr_00140 3960 3961 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00139 7514 3960 3962 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00138 3984 3986 3960 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00137 4215 3984 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00136 7514 3984 4215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00135 3962 3986 3961 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00134 3961 3988 3985 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00133 518 3081 489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00132 489 1085 518 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00131 7514 775 489 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00130 4110 4702 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00129 6549 4249 4110 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00128 5198 5214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00127 5215 6672 5198 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00126 7514 5249 5097 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00125 5097 5688 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00124 7514 5378 5097 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00123 7514 5832 4514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00122 4514 4827 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00121 7514 4511 4514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00120 7514 7224 7148 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00119 7147 7148 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00118 7514 7148 7147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00117 7514 7148 7147 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00116 7147 7148 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00115 7514 7224 7214 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00114 7213 7214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00113 7514 7214 7213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00112 7514 7214 7213 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00111 7213 7214 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00110 7514 7224 7216 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00109 7215 7216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00108 7514 7216 7215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00107 7514 7216 7215 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00106 7215 7216 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00105 7514 7224 7155 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00104 7154 7155 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00103 7514 7155 7154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00102 7514 7155 7154 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00101 7154 7155 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00100 7514 7224 7223 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00099 7222 7223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00098 7514 7223 7222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00097 7514 7223 7222 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00096 7222 7223 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00095 7514 7224 7226 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00094 7225 7226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00093 7514 7226 7225 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00092 7514 7226 7225 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00091 7225 7226 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00090 7294 7327 7313 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00089 7514 7466 7294 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00088 7295 7474 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00087 7313 7328 7295 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00086 7514 7474 7327 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00085 7328 7466 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.75U AS=0.195P AD=0.195P PS=2.02U PD=2.02U 
Mtr_00084 910 653 624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00083 624 654 910 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00082 7514 833 624 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00081 7355 7353 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00080 7354 7384 7355 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00079 3065 6340 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00078 3120 3516 3065 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00077 7514 7240 6192 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00076 6191 6192 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00075 7514 6192 6191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00074 7514 6192 6191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00073 6191 6192 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00072 880 907 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00071 908 1341 880 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00070 840 4600 839 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00069 839 1292 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00068 4368 7042 840 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00067 6764 7334 6765 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00066 6765 7383 6764 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00065 7514 6965 6765 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00064 5765 6968 5766 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00063 5766 6156 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00062 5803 7452 5765 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00061 7514 7240 6262 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00060 6261 6262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00059 7514 6262 6261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00058 7514 6262 6261 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00057 6261 6262 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00056 7514 7240 6264 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00055 6263 6264 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00054 7514 6264 6263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00053 7514 6264 6263 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00052 6263 6264 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00051 7514 7240 6200 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00050 6199 6200 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00049 7514 6200 6199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00048 7514 6200 6199 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00047 6199 6200 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00046 7514 7240 6269 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00045 6268 6269 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00044 7514 6269 6268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00043 7514 6269 6268 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00042 6268 6269 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00041 7267 7491 7266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00040 7266 7379 7267 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00039 7514 7464 7266 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00038 7514 2337 2191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00037 2191 2338 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00036 2189 2190 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00035 2191 2467 2190 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00034 2190 3837 2191 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.27U AS=0.3302P AD=0.3302P PS=3.07U PD=3.07U 
Mtr_00033 5196 5841 5195 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00032 5195 5842 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00031 5889 6333 5196 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00030 2026 2945 2025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00029 2025 2946 2026 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00028 7514 5138 2025 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00027 2099 2026 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00026 7440 7513 7186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00025 7186 7243 7440 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00024 7514 7242 7186 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.5U AS=0.39P AD=0.39P PS=3.52U PD=3.52U 
Mtr_00023 7514 7240 6270 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00022 6611 6270 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00021 7514 6270 6611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00020 7514 6270 6611 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00019 6611 6270 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00018 7514 7240 7161 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00017 7160 7161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00016 7514 7161 7160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00015 7514 7161 7160 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00014 7160 7161 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00013 7514 7240 7231 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00012 7230 7231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00011 7514 7231 7230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00010 7514 7231 7230 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00009 7230 7231 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00008 7514 7240 7233 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00007 7232 7233 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00006 7514 7233 7232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00005 7514 7233 7232 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00004 7232 7233 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00003 7514 4597 4599 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00002 4599 6576 4598 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
Mtr_00001 5459 4598 7514 7514 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.42U AS=0.3692P AD=0.3692P PS=3.37U PD=3.37U 
.ends m65_cts_r_ext

