* Spice description of o3_x2
* Spice driver version 1852071707
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:22

* INTERF i0 i1 i2 q vdd vss 


.subckt o3_x2 4 6 7 5 2 9 
* NET 2 = vdd
* NET 4 = i0
* NET 5 = q
* NET 6 = i1
* NET 7 = i2
* NET 9 = vss
Mtr_00008 5 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 2 4 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00006 1 6 3 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00005 3 7 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.55U AS=0.612P AD=0.612P PS=5.58U PD=5.58U 
Mtr_00004 5 8 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00003 8 6 9 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00002 9 4 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
Mtr_00001 9 7 8 9 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.85U AS=0.204P AD=0.204P PS=2.18U PD=2.18U 
C8 2 9 1.66309e-15
C6 4 9 1.39425e-15
C5 5 9 2.18213e-15
C4 6 9 1.38512e-15
C3 7 9 1.38512e-15
C2 8 9 2.81726e-15
C1 9 9 2.01861e-15
.ends o3_x2

