-- no model for nsnrlatch_x0
