* IOPadVdd
.subckt IOPadVdd vss vdd iovss iovdd
Xpad vdd Pad_15800W12000H
Xnclamp iovss iovdd vdd Clamp_N32N0D
Xpclamp iovss iovdd vdd Clamp_P32N0D
Xpad_guardring iovss GuardRing_N18000W13312HFF
.ends IOPadVdd
