* sff1r_x4
.subckt sff1r_x4 vss ck vdd i nrst q
Mn_ck_1 nckr ck vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ck_1 nckr ck vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_ckr_1 _net0 ckr sff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ckr_1 sff_m ckr _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_ckr_2 y ckr sff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_2 sff_s ckr _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i_1 u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i_1 u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_1 vss nckr ckr vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_nckr_1 vdd nckr ckr vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_2 sff_m nckr _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nckr_3 sff_s nckr _net8 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_2 _net7 nckr sff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_nckr_3 y nckr sff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nrst_2 _net8 nrst _net5 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nrst_1 _net4 nrst y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_nrst_1 y nrst vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nrst_2 vdd nrst _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_q_1 _net5 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_q_1 _net3 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_sffm_1 vss sff_m _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_sffm_1 vdd sff_m y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_sffs_1 vdd sff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_2 q sff_s vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_sffs_2 q sff_s vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_1 vss sff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_u_1 vdd u _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_u_1 vss u _net7 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_y_1 _net6 y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_y_1 _net2 y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends sff1r_x4
