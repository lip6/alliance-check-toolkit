* Spice description of noa22_x1
* Spice driver version 1265114907
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:05

* INTERF i0 i1 i2 nq vdd vss 


.subckt noa22_x1 5 4 3 6 1 8 
* NET 1 = vdd
* NET 3 = i2
* NET 4 = i1
* NET 5 = i0
* NET 6 = nq
* NET 8 = vss
Mtr_00006 1 3 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00005 2 4 6 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00004 6 5 2 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00003 8 3 6 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00002 6 4 7 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00001 7 5 8 8 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
C8 1 8 1.41822e-15
C7 2 8 7.32113e-16
C6 3 8 2.50714e-15
C5 4 8 1.45814e-15
C4 5 8 1.77397e-15
C3 6 8 2.07916e-15
C1 8 8 1.46971e-15
.ends noa22_x1

