* Spice description of mx2_x2
* Spice driver version 890646299
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:44

* INTERF cmd i0 i1 q vdd vss 


.subckt mx2_x2 9 5 3 4 2 10 
* NET 2 = vdd
* NET 3 = i1
* NET 4 = q
* NET 5 = i0
* NET 9 = cmd
* NET 10 = vss
Mtr_00012 4 8 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 1 11 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00010 8 9 8 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00009 2 9 11 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00008 2 3 1 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00007 8 5 2 2 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 7 5 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00005 4 8 10 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.61U AS=0.3864P AD=0.3864P PS=3.71U PD=3.71U 
Mtr_00004 8 11 7 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00003 10 9 11 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00002 6 9 8 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
Mtr_00001 10 3 6 10 sky130_fd_pr__nfet_01v8__model L=0.15U W=0.76U AS=0.1824P AD=0.1824P PS=2.01U PD=2.01U 
C10 2 10 3.3848e-15
C9 3 10 2.46609e-15
C8 4 10 2.15173e-15
C7 5 10 1.75763e-15
C4 8 10 1.74659e-15
C3 9 10 3.00631e-15
C2 10 10 2.7135e-15
C1 11 10 2.78163e-15
.ends mx2_x2

