-- no model for nor4_x0
