../rtl/reg4.vhdl