* DP8TArray_4X4
* DP8TCell
.subckt DP8TCell vdd vss wl1 wl2 bl1 bl1_n bl2 bl2_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 vdd bit bit_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 vss bit bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl1 wl1 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg1n bl1_n wl1 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2 bl2 wl2 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2n bl2_n wl2 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
.ends DP8TCell
* DP8TArray_2X1
.subckt DP8TArray_2X1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 vdd vss wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
Xinst1x0 vdd vss wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
.ends DP8TArray_2X1
* DP8TArray_2X2
.subckt DP8TArray_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TArray_2X1
Xinst0x1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X1
.ends DP8TArray_2X2
* DP8TArray_4X2
.subckt DP8TArray_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
.ends DP8TArray_4X2
* DP8TArray_4X4
.subckt DP8TArray_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X2
.ends DP8TArray_4X4
