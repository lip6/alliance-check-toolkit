* Spice description of na3_x4
* Spice driver version 1835319067
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:27:51

* INTERF i0 i1 i2 nq vdd vss 


.subckt na3_x4 7 3 6 4 1 5 
* NET 1 = vdd
* NET 3 = i1
* NET 4 = nq
* NET 5 = vss
* NET 6 = i2
* NET 7 = i0
Mtr_00012 1 2 4 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 4 2 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 1 3 10 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00009 10 6 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00008 1 7 10 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=2.63U AS=0.6312P AD=0.6312P PS=5.75U PD=5.75U 
Mtr_00007 2 10 1 1 sky130_fd_pr__pfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00006 5 2 4 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00005 4 2 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.46U AS=0.5904P AD=0.5904P PS=5.41U PD=5.41U 
Mtr_00004 8 6 9 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00003 5 3 8 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00002 2 10 5 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
Mtr_00001 9 7 10 5 sky130_fd_pr__nfet_01v8__model L=0.15U W=1.7U AS=0.408P AD=0.408P PS=3.88U PD=3.88U 
C10 1 5 2.30729e-15
C9 2 5 1.9517e-15
C8 3 5 1.74574e-15
C7 4 5 1.8477e-15
C6 5 5 2.57504e-15
C5 6 5 1.69828e-15
C4 7 5 1.7328e-15
C1 10 5 3.05063e-15
.ends na3_x4

