* BulkConn_18000WUp
* BulkConn_18000WUp
.subckt BulkConn_18000WUp vdd vss iovdd iovss

.ends BulkConn_18000WUp
