* ExampleSRAMs

* SP6TBlock_512x64_8WE
.subckt SP6TBlock_512x64_8WE clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] vss vdd q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] q[9] q[10] q[11] q[12] q[13] q[14] q[15] q[16] q[17] q[18] q[19] q[20] q[21] q[22] q[23] q[24] q[25] q[26] q[27] q[28] q[29] q[30] q[31] q[32] q[33] q[34] q[35] q[36] q[37] q[38] q[39] q[40] q[41] q[42] q[43] q[44] q[45] q[46] q[47] q[48] q[49] q[50] q[51] q[52] q[53] q[54] q[55] q[56] q[57] q[58] q[59] q[60] q[61] q[62] q[63] d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] d[8] d[9] d[10] d[11] d[12] d[13] d[14] d[15] d[16] d[17] d[18] d[19] d[20] d[21] d[22] d[23] d[24] d[25] d[26] d[27] d[28] d[29] d[30] d[31] d[32] d[33] d[34] d[35] d[36] d[37] d[38] d[39] d[40] d[41] d[42] d[43] d[44] d[45] d[46] d[47] d[48] d[49] d[50] d[51] d[52] d[53] d[54] d[55] d[56] d[57] d[58] d[59] d[60] d[61] d[62] d[63] we[0] we[1] we[2] we[3] we[4] we[5] we[6] we[7]
Xrowperiph vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] columnclk precharge_n we_en SP6TRowPeriphery_3_4_2
Xcolumnblock vss vdd columnclk precharge_n we_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] we[0] q[0] d[0] q[1] d[1] q[2] d[2] q[3] d[3] q[4] d[4] q[5] d[5] q[6] d[6] q[7] d[7] we[1] q[8] d[8] q[9] d[9] q[10] d[10] q[11] d[11] q[12] d[12] q[13] d[13] q[14] d[14] q[15] d[15] we[2] q[16] d[16] q[17] d[17] q[18] d[18] q[19] d[19] q[20] d[20] q[21] d[21] q[22] d[22] q[23] d[23] we[3] q[24] d[24] q[25] d[25] q[26] d[26] q[27] d[27] q[28] d[28] q[29] d[29] q[30] d[30] q[31] d[31] we[4] q[32] d[32] q[33] d[33] q[34] d[34] q[35] d[35] q[36] d[36] q[37] d[37] q[38] d[38] q[39] d[39] we[5] q[40] d[40] q[41] d[41] q[42] d[42] q[43] d[43] q[44] d[44] q[45] d[45] q[46] d[46] q[47] d[47] we[6] q[48] d[48] q[49] d[49] q[50] d[50] q[51] d[51] q[52] d[52] q[53] d[53] q[54] d[54] q[55] d[55] we[7] q[56] d[56] q[57] d[57] q[58] d[58] q[59] d[59] q[60] d[60] q[61] d[61] q[62] d[62] q[63] d[63] SP6TColumnBlock_128R64B4M8W
.ends SP6TBlock_512x64_8WE

* SP6TRowPeriphery_3_4_2
.subckt SP6TRowPeriphery_3_4_2 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] columnclk precharge_n we_en
Xclkgen vss vdd clk decodeclk columnclk precharge_n wl_en we_en SP6TClockGenerator
Xcoldec vss vdd decodeclk a[0] a[1] mux[0] mux[1] mux[2] mux[3] SP6TLatchedDecoder_2A2R
Xrowdec vss vdd a[2] a[3] a[4] a[5] a[6] a[7] a[8] decodeclk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] SP6TRowDecoder_3_4B
.ends SP6TRowPeriphery_3_4_2

* SP6TColumn_128R8B4M
.subckt SP6TColumn_128R8B4M vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[0] d[0] q[1] d[1] q[2] d[2] q[3] d[3] q[4] d[4] q[5] d[5] q[6] d[6] q[7] d[7] we clk we_en precharge_n mux[0] mux[1] mux[2] mux[3]
Xarray vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] SP6TArray_128X32
Xperiph vss vdd clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3] SP6TColumnPeriphery_8B4M
.ends SP6TColumn_128R8B4M

* SP6TColumnBlock_128R64B4M8W
.subckt SP6TColumnBlock_128R64B4M8W vss vdd clk precharge_n we_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] we[0] q[0] d[0] q[1] d[1] q[2] d[2] q[3] d[3] q[4] d[4] q[5] d[5] q[6] d[6] q[7] d[7] we[1] q[8] d[8] q[9] d[9] q[10] d[10] q[11] d[11] q[12] d[12] q[13] d[13] q[14] d[14] q[15] d[15] we[2] q[16] d[16] q[17] d[17] q[18] d[18] q[19] d[19] q[20] d[20] q[21] d[21] q[22] d[22] q[23] d[23] we[3] q[24] d[24] q[25] d[25] q[26] d[26] q[27] d[27] q[28] d[28] q[29] d[29] q[30] d[30] q[31] d[31] we[4] q[32] d[32] q[33] d[33] q[34] d[34] q[35] d[35] q[36] d[36] q[37] d[37] q[38] d[38] q[39] d[39] we[5] q[40] d[40] q[41] d[41] q[42] d[42] q[43] d[43] q[44] d[44] q[45] d[45] q[46] d[46] q[47] d[47] we[6] q[48] d[48] q[49] d[49] q[50] d[50] q[51] d[51] q[52] d[52] q[53] d[53] q[54] d[54] q[55] d[55] we[7] q[56] d[56] q[57] d[57] q[58] d[58] q[59] d[59] q[60] d[60] q[61] d[61] q[62] d[62] q[63] d[63]
Xcolumn[0] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[0] d[0] q[1] d[1] q[2] d[2] q[3] d[3] q[4] d[4] q[5] d[5] q[6] d[6] q[7] d[7] we[0] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[1] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[8] d[8] q[9] d[9] q[10] d[10] q[11] d[11] q[12] d[12] q[13] d[13] q[14] d[14] q[15] d[15] we[1] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[2] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[16] d[16] q[17] d[17] q[18] d[18] q[19] d[19] q[20] d[20] q[21] d[21] q[22] d[22] q[23] d[23] we[2] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[3] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[24] d[24] q[25] d[25] q[26] d[26] q[27] d[27] q[28] d[28] q[29] d[29] q[30] d[30] q[31] d[31] we[3] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[4] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[32] d[32] q[33] d[33] q[34] d[34] q[35] d[35] q[36] d[36] q[37] d[37] q[38] d[38] q[39] d[39] we[4] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[5] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[40] d[40] q[41] d[41] q[42] d[42] q[43] d[43] q[44] d[44] q[45] d[45] q[46] d[46] q[47] d[47] we[5] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[6] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[48] d[48] q[49] d[49] q[50] d[50] q[51] d[51] q[52] d[52] q[53] d[53] q[54] d[54] q[55] d[55] we[6] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
Xcolumn[7] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] q[56] d[56] q[57] d[57] q[58] d[58] q[59] d[59] q[60] d[60] q[61] d[61] q[62] d[62] q[63] d[63] we[7] clk we_en precharge_n mux[0] mux[1] mux[2] mux[3] SP6TColumn_128R8B4M
.ends SP6TColumnBlock_128R64B4M8W

* SP6TClockGenerator
.subckt SP6TClockGenerator vss vdd clk decodeclk columnclk precharge_n wl_en we_en
Xnonovl vss vdd clk firststage[0] firststage[1] firststage[2] firststage[3] firststage[4] firststage[5] firststage[6] firstpulse firststage[8] secondstage[0] secondstage[1] secondstage[2] secondstage[3] secondstage[4] secondstage[5] secondstage[6] secondpulse secondstage[8] SP6TNonOverlapClock_8S
Xdecodeclkbuf vdd vss clk decodeclk buf_x2
Xcolumnclkbuf vdd vss clk columnclk buf_x2
Xwlenbuf vdd vss firstpulse wl_en buf_x2
Xweenbuf vdd vss firstpulse we_en buf_x2
Xprechargeinv vdd vss secondpulse precharge_n inv_x2
.ends SP6TClockGenerator

* SP6TLatchedDecoder_2A2R
.subckt SP6TLatchedDecoder_2A2R vss vdd clk a[0] a[1] line[0] line[1] line[2] line[3]
Xaff[0] vdd clk vss a[0] aint[0] sff1_x4
Xaff[1] vdd clk vss a[1] aint[1] sff1_x4
Xainv[0] vdd vss aint[0] aint_n[0] inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] inv_x1
Xlinenand[0] vdd vss line_n[0] aint_n[0] aint_n[1] nand2_x0
Xlinenand[1] vdd vss line_n[1] aint[0] aint_n[1] nand2_x0
Xlinenand[2] vdd vss line_n[2] aint_n[0] aint[1] nand2_x0
Xlinenand[3] vdd vss line_n[3] aint[0] aint[1] nand2_x0
Xlineinv[0] vdd vss line_n[0] line[0] inv_x2
Xlineinv[1] vdd vss line_n[1] line[1] inv_x2
Xlineinv[2] vdd vss line_n[2] line[2] inv_x2
Xlineinv[3] vdd vss line_n[3] line[3] inv_x2
.ends SP6TLatchedDecoder_2A2R

* SP6TRowDecoder_3_4B
.subckt SP6TRowDecoder_3_4B vss vdd a[0] a[1] a[2] a[3] a[4] a[5] a[6] clk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
Xpredec vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] pd[1][0] pd[1][1] pd[1][2] pd[1][3] pd[1][4] pd[1][5] pd[1][6] pd[1][7] pd[1][8] pd[1][9] pd[1][10] pd[1][11] pd[1][12] pd[1][13] pd[1][14] pd[1][15] SP6TRowPredecoders_3_4B
Xpage[0] vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1][0] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[1] vss vdd pd[0][0] wl[8] pd[0][1] wl[9] pd[0][2] wl[10] pd[0][3] wl[11] pd[0][4] wl[12] pd[0][5] wl[13] pd[0][6] wl[14] pd[0][7] wl[15] pd[1][1] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[2] vss vdd pd[0][0] wl[16] pd[0][1] wl[17] pd[0][2] wl[18] pd[0][3] wl[19] pd[0][4] wl[20] pd[0][5] wl[21] pd[0][6] wl[22] pd[0][7] wl[23] pd[1][2] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[3] vss vdd pd[0][0] wl[24] pd[0][1] wl[25] pd[0][2] wl[26] pd[0][3] wl[27] pd[0][4] wl[28] pd[0][5] wl[29] pd[0][6] wl[30] pd[0][7] wl[31] pd[1][3] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[4] vss vdd pd[0][0] wl[32] pd[0][1] wl[33] pd[0][2] wl[34] pd[0][3] wl[35] pd[0][4] wl[36] pd[0][5] wl[37] pd[0][6] wl[38] pd[0][7] wl[39] pd[1][4] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[5] vss vdd pd[0][0] wl[40] pd[0][1] wl[41] pd[0][2] wl[42] pd[0][3] wl[43] pd[0][4] wl[44] pd[0][5] wl[45] pd[0][6] wl[46] pd[0][7] wl[47] pd[1][5] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[6] vss vdd pd[0][0] wl[48] pd[0][1] wl[49] pd[0][2] wl[50] pd[0][3] wl[51] pd[0][4] wl[52] pd[0][5] wl[53] pd[0][6] wl[54] pd[0][7] wl[55] pd[1][6] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[7] vss vdd pd[0][0] wl[56] pd[0][1] wl[57] pd[0][2] wl[58] pd[0][3] wl[59] pd[0][4] wl[60] pd[0][5] wl[61] pd[0][6] wl[62] pd[0][7] wl[63] pd[1][7] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[8] vss vdd pd[0][0] wl[64] pd[0][1] wl[65] pd[0][2] wl[66] pd[0][3] wl[67] pd[0][4] wl[68] pd[0][5] wl[69] pd[0][6] wl[70] pd[0][7] wl[71] pd[1][8] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[9] vss vdd pd[0][0] wl[72] pd[0][1] wl[73] pd[0][2] wl[74] pd[0][3] wl[75] pd[0][4] wl[76] pd[0][5] wl[77] pd[0][6] wl[78] pd[0][7] wl[79] pd[1][9] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[10] vss vdd pd[0][0] wl[80] pd[0][1] wl[81] pd[0][2] wl[82] pd[0][3] wl[83] pd[0][4] wl[84] pd[0][5] wl[85] pd[0][6] wl[86] pd[0][7] wl[87] pd[1][10] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[11] vss vdd pd[0][0] wl[88] pd[0][1] wl[89] pd[0][2] wl[90] pd[0][3] wl[91] pd[0][4] wl[92] pd[0][5] wl[93] pd[0][6] wl[94] pd[0][7] wl[95] pd[1][11] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[12] vss vdd pd[0][0] wl[96] pd[0][1] wl[97] pd[0][2] wl[98] pd[0][3] wl[99] pd[0][4] wl[100] pd[0][5] wl[101] pd[0][6] wl[102] pd[0][7] wl[103] pd[1][12] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[13] vss vdd pd[0][0] wl[104] pd[0][1] wl[105] pd[0][2] wl[106] pd[0][3] wl[107] pd[0][4] wl[108] pd[0][5] wl[109] pd[0][6] wl[110] pd[0][7] wl[111] pd[1][13] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[14] vss vdd pd[0][0] wl[112] pd[0][1] wl[113] pd[0][2] wl[114] pd[0][3] wl[115] pd[0][4] wl[116] pd[0][5] wl[117] pd[0][6] wl[118] pd[0][7] wl[119] pd[1][14] wl_en SP6TRowDecoderDriverPage_2PD8R
Xpage[15] vss vdd pd[0][0] wl[120] pd[0][1] wl[121] pd[0][2] wl[122] pd[0][3] wl[123] pd[0][4] wl[124] pd[0][5] wl[125] pd[0][6] wl[126] pd[0][7] wl[127] pd[1][15] wl_en SP6TRowDecoderDriverPage_2PD8R
.ends SP6TRowDecoder_3_4B

* SP6TNonOverlapClock_8S
.subckt SP6TNonOverlapClock_8S vss vdd clk firststage[0] firststage[1] firststage[2] firststage[3] firststage[4] firststage[5] firststage[6] firststage[7] firststage[8] secondstage[0] secondstage[1] secondstage[2] secondstage[3] secondstage[4] secondstage[5] secondstage[6] secondstage[7] secondstage[8]
Xclkinv vdd vss clk clk_n inv_x0
Xfirstnand2 vdd vss firststage[0] clk secondstage[8] nand2_x0
Xfirststage[0] vdd vss firststage[0] firststage[1] inv_x0
Xfirststage[1] vdd vss firststage[1] firststage[2] inv_x0
Xfirststage[2] vdd vss firststage[2] firststage[3] inv_x0
Xfirststage[3] vdd vss firststage[3] firststage[4] inv_x0
Xfirststage[4] vdd vss firststage[4] firststage[5] inv_x0
Xfirststage[5] vdd vss firststage[5] firststage[6] inv_x0
Xfirststage[6] vdd vss firststage[6] firststage[7] inv_x0
Xfirststage[7] vdd vss firststage[7] firststage[8] inv_x0
Xsecondnand2 vdd vss secondstage[0] clk_n firststage[8] nand2_x0
Xsecondstage[0] vdd vss secondstage[0] secondstage[1] inv_x0
Xsecondstage[1] vdd vss secondstage[1] secondstage[2] inv_x0
Xsecondstage[2] vdd vss secondstage[2] secondstage[3] inv_x0
Xsecondstage[3] vdd vss secondstage[3] secondstage[4] inv_x0
Xsecondstage[4] vdd vss secondstage[4] secondstage[5] inv_x0
Xsecondstage[5] vdd vss secondstage[5] secondstage[6] inv_x0
Xsecondstage[6] vdd vss secondstage[6] secondstage[7] inv_x0
Xsecondstage[7] vdd vss secondstage[7] secondstage[8] inv_x0
.ends SP6TNonOverlapClock_8S

* SP6TRowPredecoders_3_4B
.subckt SP6TRowPredecoders_3_4B vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] pd[1][0] pd[1][1] pd[1][2] pd[1][3] pd[1][4] pd[1][5] pd[1][6] pd[1][7] pd[1][8] pd[1][9] pd[1][10] pd[1][11] pd[1][12] pd[1][13] pd[1][14] pd[1][15]
Xaff[0] vdd clk vss a[0] aint[0] sff1_x4
Xaff[1] vdd clk vss a[1] aint[1] sff1_x4
Xaff[2] vdd clk vss a[2] aint[2] sff1_x4
Xaff[3] vdd clk vss a[3] aint[3] sff1_x4
Xaff[4] vdd clk vss a[4] aint[4] sff1_x4
Xaff[5] vdd clk vss a[5] aint[5] sff1_x4
Xaff[6] vdd clk vss a[6] aint[6] sff1_x4
Xainv[0] vdd vss aint[0] aint_n[0] inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] inv_x1
Xainv[2] vdd vss aint[2] aint_n[2] inv_x1
Xainv[3] vdd vss aint[3] aint_n[3] inv_x1
Xainv[4] vdd vss aint[4] aint_n[4] inv_x1
Xainv[5] vdd vss aint[5] aint_n[5] inv_x1
Xainv[6] vdd vss aint[6] aint_n[6] inv_x1
Xpd[0]and[0] vdd pd[0][0] vss aint_n[0] aint_n[1] aint_n[2] a3_x2
Xpd[0]and[1] vdd pd[0][1] vss aint[0] aint_n[1] aint_n[2] a3_x2
Xpd[0]and[2] vdd pd[0][2] vss aint_n[0] aint[1] aint_n[2] a3_x2
Xpd[0]and[3] vdd pd[0][3] vss aint[0] aint[1] aint_n[2] a3_x2
Xpd[0]and[4] vdd pd[0][4] vss aint_n[0] aint_n[1] aint[2] a3_x2
Xpd[0]and[5] vdd pd[0][5] vss aint[0] aint_n[1] aint[2] a3_x2
Xpd[0]and[6] vdd pd[0][6] vss aint_n[0] aint[1] aint[2] a3_x2
Xpd[0]and[7] vdd pd[0][7] vss aint[0] aint[1] aint[2] a3_x2
Xpd[1]and[0] vss pd[1][0] vdd aint_n[3] aint_n[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[1] vss pd[1][1] vdd aint[3] aint_n[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[2] vss pd[1][2] vdd aint_n[3] aint[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[3] vss pd[1][3] vdd aint[3] aint[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[4] vss pd[1][4] vdd aint_n[3] aint_n[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[5] vss pd[1][5] vdd aint[3] aint_n[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[6] vss pd[1][6] vdd aint_n[3] aint[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[7] vss pd[1][7] vdd aint[3] aint[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[8] vss pd[1][8] vdd aint_n[3] aint_n[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[9] vss pd[1][9] vdd aint[3] aint_n[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[10] vss pd[1][10] vdd aint_n[3] aint[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[11] vss pd[1][11] vdd aint[3] aint[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[12] vss pd[1][12] vdd aint_n[3] aint_n[4] aint[5] aint[6] a4_x2
Xpd[1]and[13] vss pd[1][13] vdd aint[3] aint_n[4] aint[5] aint[6] a4_x2
Xpd[1]and[14] vss pd[1][14] vdd aint_n[3] aint[4] aint[5] aint[6] a4_x2
Xpd[1]and[15] vss pd[1][15] vdd aint[3] aint[4] aint[5] aint[6] a4_x2
Xtie[0] vdd vss tie_diff_w4
Xtie[1] vdd vss tie_diff_w4
Xtie[2] vdd vss tie_diff_w4
Xtie[3] vdd vss tie_diff_w4
Xtie[4] vdd vss tie_diff_w4
Xtie[5] vdd vss tie_diff_w4
Xtie[6] vdd vss tie_diff_w4
Xtie[7] vdd vss tie_diff_w4
Xtie[8] vdd vss tie_diff_w4
Xtie[9] vdd vss tie_diff_w4
Xtie[10] vdd vss tie_diff_w4
Xtie[11] vdd vss tie_diff_w4
Xtie[12] vdd vss tie_diff_w4
Xtie[13] vdd vss tie_diff_w4
Xtie[14] vdd vss tie_diff_w4
Xtie[15] vdd vss tie_diff_w4
Xtie[16] vdd vss tie_diff_w4
Xtie[17] vdd vss tie_diff_w4
Xtie[18] vdd vss tie_diff_w4
Xtie[19] vdd vss tie_diff_w4
Xtie[20] vdd vss tie_diff_w4
Xtie[21] vdd vss tie_diff_w4
Xtie[22] vdd vss tie_diff_w4
Xtie[23] vdd vss tie_diff_w4
Xtie[24] vdd vss tie_diff_w4
Xtie[25] vdd vss tie_diff_w4
Xtie[26] vdd vss tie_diff_w4
Xtie[27] vdd vss tie_diff_w4
Xtie[28] vdd vss tie_diff_w4
Xtie[29] vdd vss tie_diff_w4
Xtie[30] vdd vss tie_diff_w4
Xtie[31] vdd vss tie_diff_w4
Xtie[32] vdd vss tie_diff_w4
Xtie[33] vdd vss tie_diff_w4
Xtie[34] vdd vss tie_diff_w4
Xtie[35] vdd vss tie_diff_w4
Xtie[36] vdd vss tie_diff_w4
Xtie[37] vdd vss tie_diff_w4
Xtie[38] vdd vss tie_diff_w4
Xtie[39] vdd vss tie_diff_w4
Xtie[40] vdd vss tie_diff_w4
Xtie[41] vdd vss tie_diff_w4
Xtie[42] vdd vss tie_diff_w4
Xtie[43] vdd vss tie_diff_w4
Xtie[44] vdd vss tie_diff_w4
Xtie[45] vdd vss tie_diff_w4
Xtie[46] vdd vss tie_diff_w4
Xtie[47] vdd vss tie_diff_w4
Xtie[48] vdd vss tie_diff_w4
Xtie[49] vdd vss tie_diff_w4
Xtie[50] vdd vss tie_diff_w4
Xtie[51] vdd vss tie_diff_w4
Xtie[52] vdd vss tie_diff_w4
Xtie[53] vdd vss tie_diff_w4
Xtie[54] vdd vss tie_diff_w4
Xtie[55] vdd vss tie_diff_w4
Xtie[56] vdd vss tie_diff_w4
Xtie[57] vdd vss tie_diff_w4
Xtie[58] vdd vss tie_diff_w4
Xtie[59] vdd vss tie_diff_w4
Xtie[60] vdd vss tie_diff_w4
Xtie[61] vdd vss tie_diff_w4
Xtie[62] vdd vss tie_diff_w4
Xtie[63] vdd vss tie_diff_w4
Xtie[64] vdd vss tie_diff_w4
Xtie[65] vdd vss tie_diff_w4
Xtie[66] vdd vss tie_diff_w4
Xtie[67] vdd vss tie_diff_w4
Xtie[68] vdd vss tie_diff_w4
Xtie[69] vdd vss tie_diff_w4
Xtie[70] vdd vss tie_diff_w4
Xtie[71] vdd vss tie_diff_w4
Xtie[72] vdd vss tie_diff_w4
Xtie[73] vdd vss tie_diff_w4
Xtie[74] vdd vss tie_diff_w4
Xtie[75] vdd vss tie_diff_w4
Xtie[76] vdd vss tie_diff_w4
Xtie[77] vdd vss tie_diff_w4
Xtie[78] vdd vss tie_diff_w4
Xtie[79] vdd vss tie_diff_w4
Xtie[80] vdd vss tie_diff_w4
Xtie[81] vdd vss tie_diff_w4
Xtie[82] vdd vss tie_diff_w4
Xtie[83] vdd vss tie_diff_w4
Xtie[84] vdd vss tie_diff_w4
Xtie[85] vdd vss tie_diff_w4
Xtie[86] vdd vss tie_diff_w4
Xtie[87] vdd vss tie_diff_w4
Xtie[88] vdd vss tie_diff_w4
Xtie[89] vdd vss tie_diff_w4
Xtie[90] vdd vss tie_diff_w4
Xtie[91] vdd vss tie_diff_w4
Xtie[92] vdd vss tie_diff_w4
Xtie[93] vdd vss tie_diff_w4
Xtie[94] vdd vss tie_diff_w4
Xtie[95] vdd vss tie_diff_w4
Xtie[96] vdd vss tie_diff_w4
Xtie[97] vdd vss tie_diff_w4
Xtie[98] vdd vss tie_diff_w4
Xtie[99] vdd vss tie_diff_w4
Xtie[100] vdd vss tie_diff_w4
Xtie[101] vdd vss tie_diff_w4
Xtie[102] vdd vss tie_diff_w4
Xtie[103] vdd vss tie_diff_w4
Xtie[104] vdd vss tie_diff_w4
Xtie[105] vdd vss tie_diff_w4
Xtie[106] vdd vss tie_diff_w4
Xtie[107] vdd vss tie_diff_w4
Xtie[108] vdd vss tie_diff_w4
.ends SP6TRowPredecoders_3_4B

* SP6TRowDecoderDriverPage_2PD8R
.subckt SP6TRowDecoderDriverPage_2PD8R vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1] wl_en
Xnand3[0] vss vdd pd[0][0] pd[1] wl_en wl_n[0] SP6TRowDecoderNand3
Xnand3[1] vss vdd pd[0][1] pd[1] wl_en wl_n[1] SP6TRowDecoderNand3
Xnand3[2] vss vdd pd[0][2] pd[1] wl_en wl_n[2] SP6TRowDecoderNand3
Xnand3[3] vss vdd pd[0][3] pd[1] wl_en wl_n[3] SP6TRowDecoderNand3
Xnand3[4] vss vdd pd[0][4] pd[1] wl_en wl_n[4] SP6TRowDecoderNand3
Xnand3[5] vss vdd pd[0][5] pd[1] wl_en wl_n[5] SP6TRowDecoderNand3
Xnand3[6] vss vdd pd[0][6] pd[1] wl_en wl_n[6] SP6TRowDecoderNand3
Xnand3[7] vss vdd pd[0][7] pd[1] wl_en wl_n[7] SP6TRowDecoderNand3
Xdrive[0] vss vdd wl_n[0] wl[0] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[1] vss vdd wl_n[1] wl[1] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[2] vss vdd wl_n[2] wl[2] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[3] vss vdd wl_n[3] wl[3] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[4] vss vdd wl_n[4] wl[4] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[5] vss vdd wl_n[5] wl[5] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[6] vss vdd wl_n[6] wl[6] SP6TWLDrive_30LN100WN30LP200WP
Xdrive[7] vss vdd wl_n[7] wl[7] SP6TWLDrive_30LN100WN30LP200WP
.ends SP6TRowDecoderDriverPage_2PD8R

* SP6TRowDecoderNand3
.subckt SP6TRowDecoderNand3 vss vdd pd[0] pd[1] wl_en wl_n
Mnmos[0] vss pd[0] int[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnmos[1] int[0] pd[1] int[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mnmos[2] int[1] wl_en wl_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.84um
Mpmos[0] vdd pd[0] wl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mpmos[1] wl_n pd[1] vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
Mpmos[2] vdd wl_en wl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.84um
.ends SP6TRowDecoderNand3

* SP6TCell
.subckt SP6TCell vdd vss wl bl bl_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 bit_n bit vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 bit_n bit vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl wl bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg2 bl_n wl bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
.ends SP6TCell

* SP6TWLDrive_30LN100WN30LP200WP
.subckt SP6TWLDrive_30LN100WN30LP200WP vss vdd wl_n wl_drive
Mnmos1 vss wl_n wl_drive vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mnmos2 wl_drive wl_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mpmos1 vdd wl_n wl_drive vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
Mpmos2 wl_drive wl_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
.ends SP6TWLDrive_30LN100WN30LP200WP

* SP6TArray_128X32
.subckt SP6TArray_128X32 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] SP6TArray_64X32
Xinst1x0 vss vdd wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] SP6TArray_64X32
.ends SP6TArray_128X32

* SP6TArray_64X32
.subckt SP6TArray_64X32 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] SP6TArray_32X32
Xinst1x0 vss vdd wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] SP6TArray_32X32
.ends SP6TArray_64X32

* SP6TArray_32X32
.subckt SP6TArray_32X32 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] SP6TArray_32X16
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] SP6TArray_32X16
.ends SP6TArray_32X32

* SP6TArray_32X16
.subckt SP6TArray_32X16 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] SP6TArray_16X16
Xinst1x0 vss vdd wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] SP6TArray_16X16
.ends SP6TArray_32X16

* SP6TArray_16X16
.subckt SP6TArray_16X16 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TArray_16X8
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] SP6TArray_16X8
.ends SP6TArray_16X16

* SP6TArray_16X8
.subckt SP6TArray_16X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TArray_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TArray_8X8
.ends SP6TArray_16X8

* SP6TArray_8X8
.subckt SP6TArray_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TArray_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TArray_8X4
.ends SP6TArray_8X8

* SP6TArray_8X4
.subckt SP6TArray_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TArray_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TArray_4X4
.ends SP6TArray_8X4

* SP6TArray_4X4
.subckt SP6TArray_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TArray_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TArray_4X2
.ends SP6TArray_4X4

* SP6TArray_4X2
.subckt SP6TArray_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TArray_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TArray_2X2
.ends SP6TArray_4X2

* SP6TArray_2X2
.subckt SP6TArray_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TArray_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TArray_2X1
.ends SP6TArray_2X2

* SP6TArray_2X1
.subckt SP6TArray_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 vdd vss wl[0] bl[0] bl_n[0] SP6TCell
Xinst1x0 vdd vss wl[1] bl[0] bl_n[0] SP6TCell
.ends SP6TArray_2X1

* SP6TColumnPeriphery_8B4M
.subckt SP6TColumnPeriphery_8B4M vss vdd clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd bl[0] bl_n[0] precharge_n SP6TPrecharge
Xprecharge[1] vdd bl[1] bl_n[1] precharge_n SP6TPrecharge
Xprecharge[2] vdd bl[2] bl_n[2] precharge_n SP6TPrecharge
Xprecharge[3] vdd bl[3] bl_n[3] precharge_n SP6TPrecharge
Xprecharge[4] vdd bl[4] bl_n[4] precharge_n SP6TPrecharge
Xprecharge[5] vdd bl[5] bl_n[5] precharge_n SP6TPrecharge
Xprecharge[6] vdd bl[6] bl_n[6] precharge_n SP6TPrecharge
Xprecharge[7] vdd bl[7] bl_n[7] precharge_n SP6TPrecharge
Xprecharge[8] vdd bl[8] bl_n[8] precharge_n SP6TPrecharge
Xprecharge[9] vdd bl[9] bl_n[9] precharge_n SP6TPrecharge
Xprecharge[10] vdd bl[10] bl_n[10] precharge_n SP6TPrecharge
Xprecharge[11] vdd bl[11] bl_n[11] precharge_n SP6TPrecharge
Xprecharge[12] vdd bl[12] bl_n[12] precharge_n SP6TPrecharge
Xprecharge[13] vdd bl[13] bl_n[13] precharge_n SP6TPrecharge
Xprecharge[14] vdd bl[14] bl_n[14] precharge_n SP6TPrecharge
Xprecharge[15] vdd bl[15] bl_n[15] precharge_n SP6TPrecharge
Xprecharge[16] vdd bl[16] bl_n[16] precharge_n SP6TPrecharge
Xprecharge[17] vdd bl[17] bl_n[17] precharge_n SP6TPrecharge
Xprecharge[18] vdd bl[18] bl_n[18] precharge_n SP6TPrecharge
Xprecharge[19] vdd bl[19] bl_n[19] precharge_n SP6TPrecharge
Xprecharge[20] vdd bl[20] bl_n[20] precharge_n SP6TPrecharge
Xprecharge[21] vdd bl[21] bl_n[21] precharge_n SP6TPrecharge
Xprecharge[22] vdd bl[22] bl_n[22] precharge_n SP6TPrecharge
Xprecharge[23] vdd bl[23] bl_n[23] precharge_n SP6TPrecharge
Xprecharge[24] vdd bl[24] bl_n[24] precharge_n SP6TPrecharge
Xprecharge[25] vdd bl[25] bl_n[25] precharge_n SP6TPrecharge
Xprecharge[26] vdd bl[26] bl_n[26] precharge_n SP6TPrecharge
Xprecharge[27] vdd bl[27] bl_n[27] precharge_n SP6TPrecharge
Xprecharge[28] vdd bl[28] bl_n[28] precharge_n SP6TPrecharge
Xprecharge[29] vdd bl[29] bl_n[29] precharge_n SP6TPrecharge
Xprecharge[30] vdd bl[30] bl_n[30] precharge_n SP6TPrecharge
Xprecharge[31] vdd bl[31] bl_n[31] precharge_n SP6TPrecharge
Xcolmux[0] bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl[0] muxbl_n[0] SP6TColMux_4C
Xcolmux[1] bl[4] bl_n[4] mux[0] bl[5] bl_n[5] mux[1] bl[6] bl_n[6] mux[2] bl[7] bl_n[7] mux[3] vss muxbl[1] muxbl_n[1] SP6TColMux_4C
Xcolmux[2] bl[8] bl_n[8] mux[0] bl[9] bl_n[9] mux[1] bl[10] bl_n[10] mux[2] bl[11] bl_n[11] mux[3] vss muxbl[2] muxbl_n[2] SP6TColMux_4C
Xcolmux[3] bl[12] bl_n[12] mux[0] bl[13] bl_n[13] mux[1] bl[14] bl_n[14] mux[2] bl[15] bl_n[15] mux[3] vss muxbl[3] muxbl_n[3] SP6TColMux_4C
Xcolmux[4] bl[16] bl_n[16] mux[0] bl[17] bl_n[17] mux[1] bl[18] bl_n[18] mux[2] bl[19] bl_n[19] mux[3] vss muxbl[4] muxbl_n[4] SP6TColMux_4C
Xcolmux[5] bl[20] bl_n[20] mux[0] bl[21] bl_n[21] mux[1] bl[22] bl_n[22] mux[2] bl[23] bl_n[23] mux[3] vss muxbl[5] muxbl_n[5] SP6TColMux_4C
Xcolmux[6] bl[24] bl_n[24] mux[0] bl[25] bl_n[25] mux[1] bl[26] bl_n[26] mux[2] bl[27] bl_n[27] mux[3] vss muxbl[6] muxbl_n[6] SP6TColMux_4C
Xcolmux[7] bl[28] bl_n[28] mux[0] bl[29] bl_n[29] mux[1] bl[30] bl_n[30] mux[2] bl[31] bl_n[31] mux[3] vss muxbl[7] muxbl_n[7] SP6TColMux_4C
Xsenseamp[0] vss vdd muxbl[0] muxbl_n[0] q[0] SP6TSenseAmp_4M
Xsenseamp[1] vss vdd muxbl[1] muxbl_n[1] q[1] SP6TSenseAmp_4M
Xsenseamp[2] vss vdd muxbl[2] muxbl_n[2] q[2] SP6TSenseAmp_4M
Xsenseamp[3] vss vdd muxbl[3] muxbl_n[3] q[3] SP6TSenseAmp_4M
Xsenseamp[4] vss vdd muxbl[4] muxbl_n[4] q[4] SP6TSenseAmp_4M
Xsenseamp[5] vss vdd muxbl[5] muxbl_n[5] q[5] SP6TSenseAmp_4M
Xsenseamp[6] vss vdd muxbl[6] muxbl_n[6] q[6] SP6TSenseAmp_4M
Xsenseamp[7] vss vdd muxbl[7] muxbl_n[7] q[7] SP6TSenseAmp_4M
Xwritedrive[0] vss vdd intclk we_n muxbl[0] muxbl_n[0] d[0] muxbl[1] muxbl_n[1] d[1] SP6TWriteDriver_4M2B
Xwritedrive[1] vss vdd intclk we_n muxbl[2] muxbl_n[2] d[2] muxbl[3] muxbl_n[3] d[3] SP6TWriteDriver_4M2B
Xwritedrive[2] vss vdd intclk we_n muxbl[4] muxbl_n[4] d[4] muxbl[5] muxbl_n[5] d[5] SP6TWriteDriver_4M2B
Xwritedrive[3] vss vdd intclk we_n muxbl[6] muxbl_n[6] d[6] muxbl[7] muxbl_n[7] d[7] SP6TWriteDriver_4M2B
Xclkwe vss vdd clk intclk we we_en we_n SP6TClockWE
.ends SP6TColumnPeriphery_8B4M

* SP6TPrecharge
.subckt SP6TPrecharge vdd bl bl_n precharge_n
Mpc1 vdd precharge_n bl vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc2 bl precharge_n bl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc3 bl_n precharge_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
.ends SP6TPrecharge

* SP6TColMux_4C
.subckt SP6TColMux_4C bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl muxbl_n
Mpgbl0 bl[0] mux[0] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln0 muxbl_n mux[0] bl_n[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl1 bl[1] mux[1] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln1 muxbl_n mux[1] bl_n[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl2 bl[2] mux[2] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln2 muxbl_n mux[2] bl_n[2] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl3 bl[3] mux[3] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln3 muxbl_n mux[3] bl_n[3] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
.ends SP6TColMux_4C

* SP6TSenseAmp_4M
.subckt SP6TSenseAmp_4M vss vdd bl bl_n q
Xlatch vss nq q vdd bl bl_n nsnrlatch_x1
Xtie vdd vss tie
.ends SP6TSenseAmp_4M

* SP6TWriteDriver_4M2B
.subckt SP6TWriteDriver_4M2B vss vdd clk we_n bl[0] bl_n[0] d[0] bl[1] bl_n[1] d[1]
Xff[0] vdd clk vss d[0] d_latched[0] sff1_x4
Xff[1] vdd clk vss d[1] d_latched[1] sff1_x4
Xnora[0] vdd vss bl_drive[0] d_latched[0] we_n nor2_x0
Xnora[1] vdd vss bl_drive[1] d_latched[1] we_n nor2_x0
Xinv[0] vdd vss d_latched[0] d_n[0] inv_x0
Xinv[1] vdd vss d_latched[1] d_n[1] inv_x0
Xnorb[0] vdd vss bln_drive[0] d_n[0] we_n nor2_x0
Xnorb[1] vdd vss bln_drive[1] d_n[1] we_n nor2_x0
Mblpd[0] vss bl_drive[0] bl[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblpd[1] vss bl_drive[1] bl[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[0] bl_n[0] bln_drive[0] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[1] bl_n[1] bln_drive[1] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
.ends SP6TWriteDriver_4M2B

* SP6TClockWE
.subckt SP6TClockWE vss vdd clkup clklow we we_en we_n
Xclkbuf vdd vss clkup clklow buf_x2
Xweff vdd clklow vss we we_latched sff1_x4
Xwenand vdd vss we_n we_en we_latched nand2_x0
.ends SP6TClockWE

* DP8TBlock_512x64_8WE
.subckt DP8TBlock_512x64_8WE clk1 clk2 a1[0] a2[0] a1[1] a2[1] a1[2] a2[2] a1[3] a2[3] a1[4] a2[4] a1[5] a2[5] a1[6] a2[6] a1[7] a2[7] a1[8] a2[8] vss vdd q1[0] q1[1] q1[2] q1[3] q1[4] q1[5] q1[6] q1[7] q1[8] q1[9] q1[10] q1[11] q1[12] q1[13] q1[14] q1[15] q1[16] q1[17] q1[18] q1[19] q1[20] q1[21] q1[22] q1[23] q1[24] q1[25] q1[26] q1[27] q1[28] q1[29] q1[30] q1[31] q1[32] q1[33] q1[34] q1[35] q1[36] q1[37] q1[38] q1[39] q1[40] q1[41] q1[42] q1[43] q1[44] q1[45] q1[46] q1[47] q1[48] q1[49] q1[50] q1[51] q1[52] q1[53] q1[54] q1[55] q1[56] q1[57] q1[58] q1[59] q1[60] q1[61] q1[62] q1[63] q2[0] q2[1] q2[2] q2[3] q2[4] q2[5] q2[6] q2[7] q2[8] q2[9] q2[10] q2[11] q2[12] q2[13] q2[14] q2[15] q2[16] q2[17] q2[18] q2[19] q2[20] q2[21] q2[22] q2[23] q2[24] q2[25] q2[26] q2[27] q2[28] q2[29] q2[30] q2[31] q2[32] q2[33] q2[34] q2[35] q2[36] q2[37] q2[38] q2[39] q2[40] q2[41] q2[42] q2[43] q2[44] q2[45] q2[46] q2[47] q2[48] q2[49] q2[50] q2[51] q2[52] q2[53] q2[54] q2[55] q2[56] q2[57] q2[58] q2[59] q2[60] q2[61] q2[62] q2[63] d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d1[6] d1[7] d1[8] d1[9] d1[10] d1[11] d1[12] d1[13] d1[14] d1[15] d1[16] d1[17] d1[18] d1[19] d1[20] d1[21] d1[22] d1[23] d1[24] d1[25] d1[26] d1[27] d1[28] d1[29] d1[30] d1[31] d1[32] d1[33] d1[34] d1[35] d1[36] d1[37] d1[38] d1[39] d1[40] d1[41] d1[42] d1[43] d1[44] d1[45] d1[46] d1[47] d1[48] d1[49] d1[50] d1[51] d1[52] d1[53] d1[54] d1[55] d1[56] d1[57] d1[58] d1[59] d1[60] d1[61] d1[62] d1[63] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5] d2[6] d2[7] d2[8] d2[9] d2[10] d2[11] d2[12] d2[13] d2[14] d2[15] d2[16] d2[17] d2[18] d2[19] d2[20] d2[21] d2[22] d2[23] d2[24] d2[25] d2[26] d2[27] d2[28] d2[29] d2[30] d2[31] d2[32] d2[33] d2[34] d2[35] d2[36] d2[37] d2[38] d2[39] d2[40] d2[41] d2[42] d2[43] d2[44] d2[45] d2[46] d2[47] d2[48] d2[49] d2[50] d2[51] d2[52] d2[53] d2[54] d2[55] d2[56] d2[57] d2[58] d2[59] d2[60] d2[61] d2[62] d2[63] we1[0] we1[1] we1[2] we1[3] we1[4] we1[5] we1[6] we1[7] we2[0] we2[1] we2[2] we2[3] we2[4] we2[5] we2[6] we2[7]
Xrowperiph1 vss vdd clk1 a1[0] a1[1] a1[2] a1[3] a1[4] a1[5] a1[6] a1[7] a1[8] wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] mux1[0] mux1[1] mux1[2] mux1[3] columnclk1 precharge1_n we_en1 DP8TRowPeriphery_3_4_2_wl1
Xrowperiph2 vss vdd clk2 a2[0] a2[1] a2[2] a2[3] a2[4] a2[5] a2[6] a2[7] a2[8] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux2[0] mux2[1] mux2[2] mux2[3] columnclk2 precharge2_n we_en2 DP8TRowPeriphery_3_4_2_wl2
Xcolumnblock vss vdd columnclk1 columnclk2 precharge1_n precharge2_n we_en1 we_en2 wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux1[0] mux1[1] mux1[2] mux1[3] mux2[0] mux2[1] mux2[2] mux2[3] we1[0] we2[0] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[1] we2[1] q1[8] q2[8] d1[8] d2[8] q1[9] q2[9] d1[9] d2[9] q1[10] q2[10] d1[10] d2[10] q1[11] q2[11] d1[11] d2[11] q1[12] q2[12] d1[12] d2[12] q1[13] q2[13] d1[13] d2[13] q1[14] q2[14] d1[14] d2[14] q1[15] q2[15] d1[15] d2[15] we1[2] we2[2] q1[16] q2[16] d1[16] d2[16] q1[17] q2[17] d1[17] d2[17] q1[18] q2[18] d1[18] d2[18] q1[19] q2[19] d1[19] d2[19] q1[20] q2[20] d1[20] d2[20] q1[21] q2[21] d1[21] d2[21] q1[22] q2[22] d1[22] d2[22] q1[23] q2[23] d1[23] d2[23] we1[3] we2[3] q1[24] q2[24] d1[24] d2[24] q1[25] q2[25] d1[25] d2[25] q1[26] q2[26] d1[26] d2[26] q1[27] q2[27] d1[27] d2[27] q1[28] q2[28] d1[28] d2[28] q1[29] q2[29] d1[29] d2[29] q1[30] q2[30] d1[30] d2[30] q1[31] q2[31] d1[31] d2[31] we1[4] we2[4] q1[32] q2[32] d1[32] d2[32] q1[33] q2[33] d1[33] d2[33] q1[34] q2[34] d1[34] d2[34] q1[35] q2[35] d1[35] d2[35] q1[36] q2[36] d1[36] d2[36] q1[37] q2[37] d1[37] d2[37] q1[38] q2[38] d1[38] d2[38] q1[39] q2[39] d1[39] d2[39] we1[5] we2[5] q1[40] q2[40] d1[40] d2[40] q1[41] q2[41] d1[41] d2[41] q1[42] q2[42] d1[42] d2[42] q1[43] q2[43] d1[43] d2[43] q1[44] q2[44] d1[44] d2[44] q1[45] q2[45] d1[45] d2[45] q1[46] q2[46] d1[46] d2[46] q1[47] q2[47] d1[47] d2[47] we1[6] we2[6] q1[48] q2[48] d1[48] d2[48] q1[49] q2[49] d1[49] d2[49] q1[50] q2[50] d1[50] d2[50] q1[51] q2[51] d1[51] d2[51] q1[52] q2[52] d1[52] d2[52] q1[53] q2[53] d1[53] d2[53] q1[54] q2[54] d1[54] d2[54] q1[55] q2[55] d1[55] d2[55] we1[7] we2[7] q1[56] q2[56] d1[56] d2[56] q1[57] q2[57] d1[57] d2[57] q1[58] q2[58] d1[58] d2[58] q1[59] q2[59] d1[59] d2[59] q1[60] q2[60] d1[60] d2[60] q1[61] q2[61] d1[61] d2[61] q1[62] q2[62] d1[62] d2[62] q1[63] q2[63] d1[63] d2[63] DP8TColumnBlock_128R64B4M8W
.ends DP8TBlock_512x64_8WE

* DP8TRowPeriphery_3_4_2_wl1
.subckt DP8TRowPeriphery_3_4_2_wl1 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] columnclk precharge_n we_en
Xclkgen vss vdd clk decodeclk columnclk precharge_n wl_en we_en DP8TClockGenerator
Xcoldec vss vdd decodeclk a[0] a[1] mux[0] mux[1] mux[2] mux[3] DP8TLatchedDecoder_2A2R
Xrowdec vss vdd a[2] a[3] a[4] a[5] a[6] a[7] a[8] decodeclk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] DP8TRowDecoder_3_4B_wl1
.ends DP8TRowPeriphery_3_4_2_wl1

* DP8TRowPeriphery_3_4_2_wl2
.subckt DP8TRowPeriphery_3_4_2_wl2 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] columnclk precharge_n we_en
Xclkgen vss vdd clk decodeclk columnclk precharge_n wl_en we_en DP8TClockGenerator
Xcoldec vss vdd decodeclk a[0] a[1] mux[0] mux[1] mux[2] mux[3] DP8TLatchedDecoder_2A2R
Xrowdec vss vdd a[2] a[3] a[4] a[5] a[6] a[7] a[8] decodeclk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] DP8TRowDecoder_3_4B_wl2
.ends DP8TRowPeriphery_3_4_2_wl2

* DP8TColumn_128R8B4M
.subckt DP8TColumn_128R8B4M vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1 clk1 we_en1 precharge1_n we2 clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3]
Xarray vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_128X32
Xperiph1 vss vdd clk1 precharge1_n we1 we_en1 q1[0] d1[0] bl1[0] bl1_n[0] bl1[1] bl1_n[1] bl1[2] bl1_n[2] bl1[3] bl1_n[3] q1[1] d1[1] bl1[4] bl1_n[4] bl1[5] bl1_n[5] bl1[6] bl1_n[6] bl1[7] bl1_n[7] q1[2] d1[2] bl1[8] bl1_n[8] bl1[9] bl1_n[9] bl1[10] bl1_n[10] bl1[11] bl1_n[11] q1[3] d1[3] bl1[12] bl1_n[12] bl1[13] bl1_n[13] bl1[14] bl1_n[14] bl1[15] bl1_n[15] q1[4] d1[4] bl1[16] bl1_n[16] bl1[17] bl1_n[17] bl1[18] bl1_n[18] bl1[19] bl1_n[19] q1[5] d1[5] bl1[20] bl1_n[20] bl1[21] bl1_n[21] bl1[22] bl1_n[22] bl1[23] bl1_n[23] q1[6] d1[6] bl1[24] bl1_n[24] bl1[25] bl1_n[25] bl1[26] bl1_n[26] bl1[27] bl1_n[27] q1[7] d1[7] bl1[28] bl1_n[28] bl1[29] bl1_n[29] bl1[30] bl1_n[30] bl1[31] bl1_n[31] mux1[0] mux1[1] mux1[2] mux1[3] DP8TColumnPeriphery_8B4M_bl1
Xperiph2 vss vdd clk2 precharge2_n we2 we_en2 q2[0] d2[0] bl2[0] bl2_n[0] bl2[1] bl2_n[1] bl2[2] bl2_n[2] bl2[3] bl2_n[3] q2[1] d2[1] bl2[4] bl2_n[4] bl2[5] bl2_n[5] bl2[6] bl2_n[6] bl2[7] bl2_n[7] q2[2] d2[2] bl2[8] bl2_n[8] bl2[9] bl2_n[9] bl2[10] bl2_n[10] bl2[11] bl2_n[11] q2[3] d2[3] bl2[12] bl2_n[12] bl2[13] bl2_n[13] bl2[14] bl2_n[14] bl2[15] bl2_n[15] q2[4] d2[4] bl2[16] bl2_n[16] bl2[17] bl2_n[17] bl2[18] bl2_n[18] bl2[19] bl2_n[19] q2[5] d2[5] bl2[20] bl2_n[20] bl2[21] bl2_n[21] bl2[22] bl2_n[22] bl2[23] bl2_n[23] q2[6] d2[6] bl2[24] bl2_n[24] bl2[25] bl2_n[25] bl2[26] bl2_n[26] bl2[27] bl2_n[27] q2[7] d2[7] bl2[28] bl2_n[28] bl2[29] bl2_n[29] bl2[30] bl2_n[30] bl2[31] bl2_n[31] mux2[0] mux2[1] mux2[2] mux2[3] DP8TColumnPeriphery_8B4M_bl2
.ends DP8TColumn_128R8B4M

* DP8TColumnBlock_128R64B4M8W
.subckt DP8TColumnBlock_128R64B4M8W vss vdd clk1 clk2 precharge1_n precharge2_n we_en1 we_en2 wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux1[0] mux1[1] mux1[2] mux1[3] mux2[0] mux2[1] mux2[2] mux2[3] we1[0] we2[0] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[1] we2[1] q1[8] q2[8] d1[8] d2[8] q1[9] q2[9] d1[9] d2[9] q1[10] q2[10] d1[10] d2[10] q1[11] q2[11] d1[11] d2[11] q1[12] q2[12] d1[12] d2[12] q1[13] q2[13] d1[13] d2[13] q1[14] q2[14] d1[14] d2[14] q1[15] q2[15] d1[15] d2[15] we1[2] we2[2] q1[16] q2[16] d1[16] d2[16] q1[17] q2[17] d1[17] d2[17] q1[18] q2[18] d1[18] d2[18] q1[19] q2[19] d1[19] d2[19] q1[20] q2[20] d1[20] d2[20] q1[21] q2[21] d1[21] d2[21] q1[22] q2[22] d1[22] d2[22] q1[23] q2[23] d1[23] d2[23] we1[3] we2[3] q1[24] q2[24] d1[24] d2[24] q1[25] q2[25] d1[25] d2[25] q1[26] q2[26] d1[26] d2[26] q1[27] q2[27] d1[27] d2[27] q1[28] q2[28] d1[28] d2[28] q1[29] q2[29] d1[29] d2[29] q1[30] q2[30] d1[30] d2[30] q1[31] q2[31] d1[31] d2[31] we1[4] we2[4] q1[32] q2[32] d1[32] d2[32] q1[33] q2[33] d1[33] d2[33] q1[34] q2[34] d1[34] d2[34] q1[35] q2[35] d1[35] d2[35] q1[36] q2[36] d1[36] d2[36] q1[37] q2[37] d1[37] d2[37] q1[38] q2[38] d1[38] d2[38] q1[39] q2[39] d1[39] d2[39] we1[5] we2[5] q1[40] q2[40] d1[40] d2[40] q1[41] q2[41] d1[41] d2[41] q1[42] q2[42] d1[42] d2[42] q1[43] q2[43] d1[43] d2[43] q1[44] q2[44] d1[44] d2[44] q1[45] q2[45] d1[45] d2[45] q1[46] q2[46] d1[46] d2[46] q1[47] q2[47] d1[47] d2[47] we1[6] we2[6] q1[48] q2[48] d1[48] d2[48] q1[49] q2[49] d1[49] d2[49] q1[50] q2[50] d1[50] d2[50] q1[51] q2[51] d1[51] d2[51] q1[52] q2[52] d1[52] d2[52] q1[53] q2[53] d1[53] d2[53] q1[54] q2[54] d1[54] d2[54] q1[55] q2[55] d1[55] d2[55] we1[7] we2[7] q1[56] q2[56] d1[56] d2[56] q1[57] q2[57] d1[57] d2[57] q1[58] q2[58] d1[58] d2[58] q1[59] q2[59] d1[59] d2[59] q1[60] q2[60] d1[60] d2[60] q1[61] q2[61] d1[61] d2[61] q1[62] q2[62] d1[62] d2[62] q1[63] q2[63] d1[63] d2[63]
Xcolumn[0] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[0] clk1 we_en1 precharge1_n we2[0] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[1] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[8] q2[8] d1[8] d2[8] q1[9] q2[9] d1[9] d2[9] q1[10] q2[10] d1[10] d2[10] q1[11] q2[11] d1[11] d2[11] q1[12] q2[12] d1[12] d2[12] q1[13] q2[13] d1[13] d2[13] q1[14] q2[14] d1[14] d2[14] q1[15] q2[15] d1[15] d2[15] we1[1] clk1 we_en1 precharge1_n we2[1] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[2] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[16] q2[16] d1[16] d2[16] q1[17] q2[17] d1[17] d2[17] q1[18] q2[18] d1[18] d2[18] q1[19] q2[19] d1[19] d2[19] q1[20] q2[20] d1[20] d2[20] q1[21] q2[21] d1[21] d2[21] q1[22] q2[22] d1[22] d2[22] q1[23] q2[23] d1[23] d2[23] we1[2] clk1 we_en1 precharge1_n we2[2] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[3] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[24] q2[24] d1[24] d2[24] q1[25] q2[25] d1[25] d2[25] q1[26] q2[26] d1[26] d2[26] q1[27] q2[27] d1[27] d2[27] q1[28] q2[28] d1[28] d2[28] q1[29] q2[29] d1[29] d2[29] q1[30] q2[30] d1[30] d2[30] q1[31] q2[31] d1[31] d2[31] we1[3] clk1 we_en1 precharge1_n we2[3] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[4] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[32] q2[32] d1[32] d2[32] q1[33] q2[33] d1[33] d2[33] q1[34] q2[34] d1[34] d2[34] q1[35] q2[35] d1[35] d2[35] q1[36] q2[36] d1[36] d2[36] q1[37] q2[37] d1[37] d2[37] q1[38] q2[38] d1[38] d2[38] q1[39] q2[39] d1[39] d2[39] we1[4] clk1 we_en1 precharge1_n we2[4] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[5] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[40] q2[40] d1[40] d2[40] q1[41] q2[41] d1[41] d2[41] q1[42] q2[42] d1[42] d2[42] q1[43] q2[43] d1[43] d2[43] q1[44] q2[44] d1[44] d2[44] q1[45] q2[45] d1[45] d2[45] q1[46] q2[46] d1[46] d2[46] q1[47] q2[47] d1[47] d2[47] we1[5] clk1 we_en1 precharge1_n we2[5] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[6] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[48] q2[48] d1[48] d2[48] q1[49] q2[49] d1[49] d2[49] q1[50] q2[50] d1[50] d2[50] q1[51] q2[51] d1[51] d2[51] q1[52] q2[52] d1[52] d2[52] q1[53] q2[53] d1[53] d2[53] q1[54] q2[54] d1[54] d2[54] q1[55] q2[55] d1[55] d2[55] we1[6] clk1 we_en1 precharge1_n we2[6] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
Xcolumn[7] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[56] q2[56] d1[56] d2[56] q1[57] q2[57] d1[57] d2[57] q1[58] q2[58] d1[58] d2[58] q1[59] q2[59] d1[59] d2[59] q1[60] q2[60] d1[60] d2[60] q1[61] q2[61] d1[61] d2[61] q1[62] q2[62] d1[62] d2[62] q1[63] q2[63] d1[63] d2[63] we1[7] clk1 we_en1 precharge1_n we2[7] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
.ends DP8TColumnBlock_128R64B4M8W

* DP8TClockGenerator
.subckt DP8TClockGenerator vss vdd clk decodeclk columnclk precharge_n wl_en we_en
Xnonovl vss vdd clk firststage[0] firststage[1] firststage[2] firststage[3] firststage[4] firststage[5] firststage[6] firstpulse firststage[8] secondstage[0] secondstage[1] secondstage[2] secondstage[3] secondstage[4] secondstage[5] secondstage[6] secondpulse secondstage[8] DP8TNonOverlapClock_8S
Xdecodeclkbuf vdd vss clk decodeclk buf_x2
Xcolumnclkbuf vdd vss clk columnclk buf_x2
Xwlenbuf vdd vss firstpulse wl_en buf_x2
Xweenbuf vdd vss firstpulse we_en buf_x2
Xprechargeinv vdd vss secondpulse precharge_n inv_x2
.ends DP8TClockGenerator

* DP8TLatchedDecoder_2A2R
.subckt DP8TLatchedDecoder_2A2R vss vdd clk a[0] a[1] line[0] line[1] line[2] line[3]
Xaff[0] vdd clk vss a[0] aint[0] sff1_x4
Xaff[1] vdd clk vss a[1] aint[1] sff1_x4
Xainv[0] vdd vss aint[0] aint_n[0] inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] inv_x1
Xlinenand[0] vdd vss line_n[0] aint_n[0] aint_n[1] nand2_x0
Xlinenand[1] vdd vss line_n[1] aint[0] aint_n[1] nand2_x0
Xlinenand[2] vdd vss line_n[2] aint_n[0] aint[1] nand2_x0
Xlinenand[3] vdd vss line_n[3] aint[0] aint[1] nand2_x0
Xlineinv[0] vdd vss line_n[0] line[0] inv_x2
Xlineinv[1] vdd vss line_n[1] line[1] inv_x2
Xlineinv[2] vdd vss line_n[2] line[2] inv_x2
Xlineinv[3] vdd vss line_n[3] line[3] inv_x2
.ends DP8TLatchedDecoder_2A2R

* DP8TRowDecoder_3_4B_wl1
.subckt DP8TRowDecoder_3_4B_wl1 vss vdd a[0] a[1] a[2] a[3] a[4] a[5] a[6] clk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
Xpredec vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] pd[1][0] pd[1][1] pd[1][2] pd[1][3] pd[1][4] pd[1][5] pd[1][6] pd[1][7] pd[1][8] pd[1][9] pd[1][10] pd[1][11] pd[1][12] pd[1][13] pd[1][14] pd[1][15] DP8TRowPredecoders_3_4B
Xpage[0] vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1][0] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[1] vss vdd pd[0][0] wl[8] pd[0][1] wl[9] pd[0][2] wl[10] pd[0][3] wl[11] pd[0][4] wl[12] pd[0][5] wl[13] pd[0][6] wl[14] pd[0][7] wl[15] pd[1][1] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[2] vss vdd pd[0][0] wl[16] pd[0][1] wl[17] pd[0][2] wl[18] pd[0][3] wl[19] pd[0][4] wl[20] pd[0][5] wl[21] pd[0][6] wl[22] pd[0][7] wl[23] pd[1][2] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[3] vss vdd pd[0][0] wl[24] pd[0][1] wl[25] pd[0][2] wl[26] pd[0][3] wl[27] pd[0][4] wl[28] pd[0][5] wl[29] pd[0][6] wl[30] pd[0][7] wl[31] pd[1][3] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[4] vss vdd pd[0][0] wl[32] pd[0][1] wl[33] pd[0][2] wl[34] pd[0][3] wl[35] pd[0][4] wl[36] pd[0][5] wl[37] pd[0][6] wl[38] pd[0][7] wl[39] pd[1][4] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[5] vss vdd pd[0][0] wl[40] pd[0][1] wl[41] pd[0][2] wl[42] pd[0][3] wl[43] pd[0][4] wl[44] pd[0][5] wl[45] pd[0][6] wl[46] pd[0][7] wl[47] pd[1][5] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[6] vss vdd pd[0][0] wl[48] pd[0][1] wl[49] pd[0][2] wl[50] pd[0][3] wl[51] pd[0][4] wl[52] pd[0][5] wl[53] pd[0][6] wl[54] pd[0][7] wl[55] pd[1][6] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[7] vss vdd pd[0][0] wl[56] pd[0][1] wl[57] pd[0][2] wl[58] pd[0][3] wl[59] pd[0][4] wl[60] pd[0][5] wl[61] pd[0][6] wl[62] pd[0][7] wl[63] pd[1][7] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[8] vss vdd pd[0][0] wl[64] pd[0][1] wl[65] pd[0][2] wl[66] pd[0][3] wl[67] pd[0][4] wl[68] pd[0][5] wl[69] pd[0][6] wl[70] pd[0][7] wl[71] pd[1][8] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[9] vss vdd pd[0][0] wl[72] pd[0][1] wl[73] pd[0][2] wl[74] pd[0][3] wl[75] pd[0][4] wl[76] pd[0][5] wl[77] pd[0][6] wl[78] pd[0][7] wl[79] pd[1][9] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[10] vss vdd pd[0][0] wl[80] pd[0][1] wl[81] pd[0][2] wl[82] pd[0][3] wl[83] pd[0][4] wl[84] pd[0][5] wl[85] pd[0][6] wl[86] pd[0][7] wl[87] pd[1][10] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[11] vss vdd pd[0][0] wl[88] pd[0][1] wl[89] pd[0][2] wl[90] pd[0][3] wl[91] pd[0][4] wl[92] pd[0][5] wl[93] pd[0][6] wl[94] pd[0][7] wl[95] pd[1][11] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[12] vss vdd pd[0][0] wl[96] pd[0][1] wl[97] pd[0][2] wl[98] pd[0][3] wl[99] pd[0][4] wl[100] pd[0][5] wl[101] pd[0][6] wl[102] pd[0][7] wl[103] pd[1][12] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[13] vss vdd pd[0][0] wl[104] pd[0][1] wl[105] pd[0][2] wl[106] pd[0][3] wl[107] pd[0][4] wl[108] pd[0][5] wl[109] pd[0][6] wl[110] pd[0][7] wl[111] pd[1][13] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[14] vss vdd pd[0][0] wl[112] pd[0][1] wl[113] pd[0][2] wl[114] pd[0][3] wl[115] pd[0][4] wl[116] pd[0][5] wl[117] pd[0][6] wl[118] pd[0][7] wl[119] pd[1][14] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[15] vss vdd pd[0][0] wl[120] pd[0][1] wl[121] pd[0][2] wl[122] pd[0][3] wl[123] pd[0][4] wl[124] pd[0][5] wl[125] pd[0][6] wl[126] pd[0][7] wl[127] pd[1][15] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
.ends DP8TRowDecoder_3_4B_wl1

* DP8TNonOverlapClock_8S
.subckt DP8TNonOverlapClock_8S vss vdd clk firststage[0] firststage[1] firststage[2] firststage[3] firststage[4] firststage[5] firststage[6] firststage[7] firststage[8] secondstage[0] secondstage[1] secondstage[2] secondstage[3] secondstage[4] secondstage[5] secondstage[6] secondstage[7] secondstage[8]
Xclkinv vdd vss clk clk_n inv_x0
Xfirstnand2 vdd vss firststage[0] clk secondstage[8] nand2_x0
Xfirststage[0] vdd vss firststage[0] firststage[1] inv_x0
Xfirststage[1] vdd vss firststage[1] firststage[2] inv_x0
Xfirststage[2] vdd vss firststage[2] firststage[3] inv_x0
Xfirststage[3] vdd vss firststage[3] firststage[4] inv_x0
Xfirststage[4] vdd vss firststage[4] firststage[5] inv_x0
Xfirststage[5] vdd vss firststage[5] firststage[6] inv_x0
Xfirststage[6] vdd vss firststage[6] firststage[7] inv_x0
Xfirststage[7] vdd vss firststage[7] firststage[8] inv_x0
Xsecondnand2 vdd vss secondstage[0] clk_n firststage[8] nand2_x0
Xsecondstage[0] vdd vss secondstage[0] secondstage[1] inv_x0
Xsecondstage[1] vdd vss secondstage[1] secondstage[2] inv_x0
Xsecondstage[2] vdd vss secondstage[2] secondstage[3] inv_x0
Xsecondstage[3] vdd vss secondstage[3] secondstage[4] inv_x0
Xsecondstage[4] vdd vss secondstage[4] secondstage[5] inv_x0
Xsecondstage[5] vdd vss secondstage[5] secondstage[6] inv_x0
Xsecondstage[6] vdd vss secondstage[6] secondstage[7] inv_x0
Xsecondstage[7] vdd vss secondstage[7] secondstage[8] inv_x0
.ends DP8TNonOverlapClock_8S

* DP8TRowPredecoders_3_4B
.subckt DP8TRowPredecoders_3_4B vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] pd[1][0] pd[1][1] pd[1][2] pd[1][3] pd[1][4] pd[1][5] pd[1][6] pd[1][7] pd[1][8] pd[1][9] pd[1][10] pd[1][11] pd[1][12] pd[1][13] pd[1][14] pd[1][15]
Xaff[0] vdd clk vss a[0] aint[0] sff1_x4
Xaff[1] vdd clk vss a[1] aint[1] sff1_x4
Xaff[2] vdd clk vss a[2] aint[2] sff1_x4
Xaff[3] vdd clk vss a[3] aint[3] sff1_x4
Xaff[4] vdd clk vss a[4] aint[4] sff1_x4
Xaff[5] vdd clk vss a[5] aint[5] sff1_x4
Xaff[6] vdd clk vss a[6] aint[6] sff1_x4
Xainv[0] vdd vss aint[0] aint_n[0] inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] inv_x1
Xainv[2] vdd vss aint[2] aint_n[2] inv_x1
Xainv[3] vdd vss aint[3] aint_n[3] inv_x1
Xainv[4] vdd vss aint[4] aint_n[4] inv_x1
Xainv[5] vdd vss aint[5] aint_n[5] inv_x1
Xainv[6] vdd vss aint[6] aint_n[6] inv_x1
Xpd[0]and[0] vdd pd[0][0] vss aint_n[0] aint_n[1] aint_n[2] a3_x2
Xpd[0]and[1] vdd pd[0][1] vss aint[0] aint_n[1] aint_n[2] a3_x2
Xpd[0]and[2] vdd pd[0][2] vss aint_n[0] aint[1] aint_n[2] a3_x2
Xpd[0]and[3] vdd pd[0][3] vss aint[0] aint[1] aint_n[2] a3_x2
Xpd[0]and[4] vdd pd[0][4] vss aint_n[0] aint_n[1] aint[2] a3_x2
Xpd[0]and[5] vdd pd[0][5] vss aint[0] aint_n[1] aint[2] a3_x2
Xpd[0]and[6] vdd pd[0][6] vss aint_n[0] aint[1] aint[2] a3_x2
Xpd[0]and[7] vdd pd[0][7] vss aint[0] aint[1] aint[2] a3_x2
Xpd[1]and[0] vss pd[1][0] vdd aint_n[3] aint_n[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[1] vss pd[1][1] vdd aint[3] aint_n[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[2] vss pd[1][2] vdd aint_n[3] aint[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[3] vss pd[1][3] vdd aint[3] aint[4] aint_n[5] aint_n[6] a4_x2
Xpd[1]and[4] vss pd[1][4] vdd aint_n[3] aint_n[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[5] vss pd[1][5] vdd aint[3] aint_n[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[6] vss pd[1][6] vdd aint_n[3] aint[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[7] vss pd[1][7] vdd aint[3] aint[4] aint[5] aint_n[6] a4_x2
Xpd[1]and[8] vss pd[1][8] vdd aint_n[3] aint_n[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[9] vss pd[1][9] vdd aint[3] aint_n[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[10] vss pd[1][10] vdd aint_n[3] aint[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[11] vss pd[1][11] vdd aint[3] aint[4] aint_n[5] aint[6] a4_x2
Xpd[1]and[12] vss pd[1][12] vdd aint_n[3] aint_n[4] aint[5] aint[6] a4_x2
Xpd[1]and[13] vss pd[1][13] vdd aint[3] aint_n[4] aint[5] aint[6] a4_x2
Xpd[1]and[14] vss pd[1][14] vdd aint_n[3] aint[4] aint[5] aint[6] a4_x2
Xpd[1]and[15] vss pd[1][15] vdd aint[3] aint[4] aint[5] aint[6] a4_x2
Xtie[0] vdd vss tie_diff_w4
Xtie[1] vdd vss tie_diff_w4
Xtie[2] vdd vss tie_diff_w4
Xtie[3] vdd vss tie_diff_w4
Xtie[4] vdd vss tie_diff_w4
Xtie[5] vdd vss tie_diff_w4
Xtie[6] vdd vss tie_diff_w4
Xtie[7] vdd vss tie_diff_w4
Xtie[8] vdd vss tie_diff_w4
Xtie[9] vdd vss tie_diff_w4
Xtie[10] vdd vss tie_diff_w4
Xtie[11] vdd vss tie_diff_w4
Xtie[12] vdd vss tie_diff_w4
Xtie[13] vdd vss tie_diff_w4
Xtie[14] vdd vss tie_diff_w4
Xtie[15] vdd vss tie_diff_w4
Xtie[16] vdd vss tie_diff_w4
Xtie[17] vdd vss tie_diff_w4
Xtie[18] vdd vss tie_diff_w4
Xtie[19] vdd vss tie_diff_w4
Xtie[20] vdd vss tie_diff_w4
Xtie[21] vdd vss tie_diff_w4
Xtie[22] vdd vss tie_diff_w4
Xtie[23] vdd vss tie_diff_w4
Xtie[24] vdd vss tie_diff_w4
Xtie[25] vdd vss tie_diff_w4
Xtie[26] vdd vss tie_diff_w4
Xtie[27] vdd vss tie_diff_w4
Xtie[28] vdd vss tie_diff_w4
Xtie[29] vdd vss tie_diff_w4
Xtie[30] vdd vss tie_diff_w4
Xtie[31] vdd vss tie_diff_w4
Xtie[32] vdd vss tie_diff_w4
Xtie[33] vdd vss tie_diff_w4
Xtie[34] vdd vss tie_diff_w4
Xtie[35] vdd vss tie_diff_w4
Xtie[36] vdd vss tie_diff_w4
Xtie[37] vdd vss tie_diff_w4
Xtie[38] vdd vss tie_diff_w4
Xtie[39] vdd vss tie_diff_w4
Xtie[40] vdd vss tie_diff_w4
Xtie[41] vdd vss tie_diff_w4
Xtie[42] vdd vss tie_diff_w4
Xtie[43] vdd vss tie_diff_w4
Xtie[44] vdd vss tie_diff_w4
Xtie[45] vdd vss tie_diff_w4
Xtie[46] vdd vss tie_diff_w4
Xtie[47] vdd vss tie_diff_w4
Xtie[48] vdd vss tie_diff_w4
Xtie[49] vdd vss tie_diff_w4
Xtie[50] vdd vss tie_diff_w4
Xtie[51] vdd vss tie_diff_w4
Xtie[52] vdd vss tie_diff_w4
Xtie[53] vdd vss tie_diff_w4
Xtie[54] vdd vss tie_diff_w4
Xtie[55] vdd vss tie_diff_w4
Xtie[56] vdd vss tie_diff_w4
Xtie[57] vdd vss tie_diff_w4
Xtie[58] vdd vss tie_diff_w4
Xtie[59] vdd vss tie_diff_w4
Xtie[60] vdd vss tie_diff_w4
Xtie[61] vdd vss tie_diff_w4
Xtie[62] vdd vss tie_diff_w4
Xtie[63] vdd vss tie_diff_w4
Xtie[64] vdd vss tie_diff_w4
Xtie[65] vdd vss tie_diff_w4
Xtie[66] vdd vss tie_diff_w4
Xtie[67] vdd vss tie_diff_w4
Xtie[68] vdd vss tie_diff_w4
Xtie[69] vdd vss tie_diff_w4
Xtie[70] vdd vss tie_diff_w4
Xtie[71] vdd vss tie_diff_w4
Xtie[72] vdd vss tie_diff_w4
Xtie[73] vdd vss tie_diff_w4
Xtie[74] vdd vss tie_diff_w4
Xtie[75] vdd vss tie_diff_w4
Xtie[76] vdd vss tie_diff_w4
Xtie[77] vdd vss tie_diff_w4
Xtie[78] vdd vss tie_diff_w4
Xtie[79] vdd vss tie_diff_w4
Xtie[80] vdd vss tie_diff_w4
Xtie[81] vdd vss tie_diff_w4
Xtie[82] vdd vss tie_diff_w4
Xtie[83] vdd vss tie_diff_w4
.ends DP8TRowPredecoders_3_4B

* DP8TRowDecoderDriverPage_2PD8R_wl1
.subckt DP8TRowDecoderDriverPage_2PD8R_wl1 vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1] wl_en
Xnand3[0] vss vdd pd[0][0] pd[1] wl_en wl_n[0] DP8TRowDecoderNand3
Xnand3[1] vss vdd pd[0][1] pd[1] wl_en wl_n[1] DP8TRowDecoderNand3
Xnand3[2] vss vdd pd[0][2] pd[1] wl_en wl_n[2] DP8TRowDecoderNand3
Xnand3[3] vss vdd pd[0][3] pd[1] wl_en wl_n[3] DP8TRowDecoderNand3
Xnand3[4] vss vdd pd[0][4] pd[1] wl_en wl_n[4] DP8TRowDecoderNand3
Xnand3[5] vss vdd pd[0][5] pd[1] wl_en wl_n[5] DP8TRowDecoderNand3
Xnand3[6] vss vdd pd[0][6] pd[1] wl_en wl_n[6] DP8TRowDecoderNand3
Xnand3[7] vss vdd pd[0][7] pd[1] wl_en wl_n[7] DP8TRowDecoderNand3
Xdrive[0] vss vdd wl_n[0] wl[0] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[1] vss vdd wl_n[1] wl[1] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[2] vss vdd wl_n[2] wl[2] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[3] vss vdd wl_n[3] wl[3] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[4] vss vdd wl_n[4] wl[4] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[5] vss vdd wl_n[5] wl[5] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[6] vss vdd wl_n[6] wl[6] DP8TWLDrive_30LN100WN30LP200WP_wl1
Xdrive[7] vss vdd wl_n[7] wl[7] DP8TWLDrive_30LN100WN30LP200WP_wl1
.ends DP8TRowDecoderDriverPage_2PD8R_wl1

* DP8TRowDecoderNand3
.subckt DP8TRowDecoderNand3 vss vdd pd[0] pd[1] wl_en wl_n
Mnmos[0] vss pd[0] int[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.65um
Mnmos[1] int[0] pd[1] int[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.65um
Mnmos[2] int[1] wl_en wl_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.65um
Mpmos[0] vdd pd[0] wl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.65um
Mpmos[1] wl_n pd[1] vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.65um
Mpmos[2] vdd wl_en wl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.65um
.ends DP8TRowDecoderNand3

* DP8TCell
.subckt DP8TCell vdd vss wl1 wl2 bl1 bl1_n bl2 bl2_n
Mpu1 vdd bit_n bit vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpu2 vdd bit bit_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpd1 vss bit_n bit vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpd2 vss bit bit_n vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.36um
Mpg1 bl1 wl1 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg1n bl1_n wl1 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2 bl2 wl2 bit vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
Mpg2n bl2_n wl2 bit_n vss sky130_fd_pr__nfet_01v8__model l=0.17um w=0.36um
.ends DP8TCell

* DP8TWLDrive_30LN100WN30LP200WP_wl1
.subckt DP8TWLDrive_30LN100WN30LP200WP_wl1 vss vdd wl_n wl_drive
Mnmos1 vss wl_n wl_drive vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mnmos2 wl_drive wl_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mpmos1 vdd wl_n wl_drive vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
Mpmos2 wl_drive wl_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
.ends DP8TWLDrive_30LN100WN30LP200WP_wl1

* DP8TRowDecoder_3_4B_wl2
.subckt DP8TRowDecoder_3_4B_wl2 vss vdd a[0] a[1] a[2] a[3] a[4] a[5] a[6] clk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
Xpredec vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] pd[1][0] pd[1][1] pd[1][2] pd[1][3] pd[1][4] pd[1][5] pd[1][6] pd[1][7] pd[1][8] pd[1][9] pd[1][10] pd[1][11] pd[1][12] pd[1][13] pd[1][14] pd[1][15] DP8TRowPredecoders_3_4B
Xpage[0] vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1][0] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[1] vss vdd pd[0][0] wl[8] pd[0][1] wl[9] pd[0][2] wl[10] pd[0][3] wl[11] pd[0][4] wl[12] pd[0][5] wl[13] pd[0][6] wl[14] pd[0][7] wl[15] pd[1][1] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[2] vss vdd pd[0][0] wl[16] pd[0][1] wl[17] pd[0][2] wl[18] pd[0][3] wl[19] pd[0][4] wl[20] pd[0][5] wl[21] pd[0][6] wl[22] pd[0][7] wl[23] pd[1][2] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[3] vss vdd pd[0][0] wl[24] pd[0][1] wl[25] pd[0][2] wl[26] pd[0][3] wl[27] pd[0][4] wl[28] pd[0][5] wl[29] pd[0][6] wl[30] pd[0][7] wl[31] pd[1][3] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[4] vss vdd pd[0][0] wl[32] pd[0][1] wl[33] pd[0][2] wl[34] pd[0][3] wl[35] pd[0][4] wl[36] pd[0][5] wl[37] pd[0][6] wl[38] pd[0][7] wl[39] pd[1][4] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[5] vss vdd pd[0][0] wl[40] pd[0][1] wl[41] pd[0][2] wl[42] pd[0][3] wl[43] pd[0][4] wl[44] pd[0][5] wl[45] pd[0][6] wl[46] pd[0][7] wl[47] pd[1][5] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[6] vss vdd pd[0][0] wl[48] pd[0][1] wl[49] pd[0][2] wl[50] pd[0][3] wl[51] pd[0][4] wl[52] pd[0][5] wl[53] pd[0][6] wl[54] pd[0][7] wl[55] pd[1][6] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[7] vss vdd pd[0][0] wl[56] pd[0][1] wl[57] pd[0][2] wl[58] pd[0][3] wl[59] pd[0][4] wl[60] pd[0][5] wl[61] pd[0][6] wl[62] pd[0][7] wl[63] pd[1][7] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[8] vss vdd pd[0][0] wl[64] pd[0][1] wl[65] pd[0][2] wl[66] pd[0][3] wl[67] pd[0][4] wl[68] pd[0][5] wl[69] pd[0][6] wl[70] pd[0][7] wl[71] pd[1][8] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[9] vss vdd pd[0][0] wl[72] pd[0][1] wl[73] pd[0][2] wl[74] pd[0][3] wl[75] pd[0][4] wl[76] pd[0][5] wl[77] pd[0][6] wl[78] pd[0][7] wl[79] pd[1][9] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[10] vss vdd pd[0][0] wl[80] pd[0][1] wl[81] pd[0][2] wl[82] pd[0][3] wl[83] pd[0][4] wl[84] pd[0][5] wl[85] pd[0][6] wl[86] pd[0][7] wl[87] pd[1][10] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[11] vss vdd pd[0][0] wl[88] pd[0][1] wl[89] pd[0][2] wl[90] pd[0][3] wl[91] pd[0][4] wl[92] pd[0][5] wl[93] pd[0][6] wl[94] pd[0][7] wl[95] pd[1][11] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[12] vss vdd pd[0][0] wl[96] pd[0][1] wl[97] pd[0][2] wl[98] pd[0][3] wl[99] pd[0][4] wl[100] pd[0][5] wl[101] pd[0][6] wl[102] pd[0][7] wl[103] pd[1][12] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[13] vss vdd pd[0][0] wl[104] pd[0][1] wl[105] pd[0][2] wl[106] pd[0][3] wl[107] pd[0][4] wl[108] pd[0][5] wl[109] pd[0][6] wl[110] pd[0][7] wl[111] pd[1][13] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[14] vss vdd pd[0][0] wl[112] pd[0][1] wl[113] pd[0][2] wl[114] pd[0][3] wl[115] pd[0][4] wl[116] pd[0][5] wl[117] pd[0][6] wl[118] pd[0][7] wl[119] pd[1][14] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[15] vss vdd pd[0][0] wl[120] pd[0][1] wl[121] pd[0][2] wl[122] pd[0][3] wl[123] pd[0][4] wl[124] pd[0][5] wl[125] pd[0][6] wl[126] pd[0][7] wl[127] pd[1][15] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
.ends DP8TRowDecoder_3_4B_wl2

* DP8TRowDecoderDriverPage_2PD8R_wl2
.subckt DP8TRowDecoderDriverPage_2PD8R_wl2 vss vdd pd[0][0] wl[0] pd[0][1] wl[1] pd[0][2] wl[2] pd[0][3] wl[3] pd[0][4] wl[4] pd[0][5] wl[5] pd[0][6] wl[6] pd[0][7] wl[7] pd[1] wl_en
Xnand3[0] vss vdd pd[0][0] pd[1] wl_en wl_n[0] DP8TRowDecoderNand3
Xnand3[1] vss vdd pd[0][1] pd[1] wl_en wl_n[1] DP8TRowDecoderNand3
Xnand3[2] vss vdd pd[0][2] pd[1] wl_en wl_n[2] DP8TRowDecoderNand3
Xnand3[3] vss vdd pd[0][3] pd[1] wl_en wl_n[3] DP8TRowDecoderNand3
Xnand3[4] vss vdd pd[0][4] pd[1] wl_en wl_n[4] DP8TRowDecoderNand3
Xnand3[5] vss vdd pd[0][5] pd[1] wl_en wl_n[5] DP8TRowDecoderNand3
Xnand3[6] vss vdd pd[0][6] pd[1] wl_en wl_n[6] DP8TRowDecoderNand3
Xnand3[7] vss vdd pd[0][7] pd[1] wl_en wl_n[7] DP8TRowDecoderNand3
Xdrive[0] vss vdd wl_n[0] wl[0] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[1] vss vdd wl_n[1] wl[1] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[2] vss vdd wl_n[2] wl[2] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[3] vss vdd wl_n[3] wl[3] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[4] vss vdd wl_n[4] wl[4] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[5] vss vdd wl_n[5] wl[5] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[6] vss vdd wl_n[6] wl[6] DP8TWLDrive_30LN100WN30LP200WP_wl2
Xdrive[7] vss vdd wl_n[7] wl[7] DP8TWLDrive_30LN100WN30LP200WP_wl2
.ends DP8TRowDecoderDriverPage_2PD8R_wl2

* DP8TWLDrive_30LN100WN30LP200WP_wl2
.subckt DP8TWLDrive_30LN100WN30LP200WP_wl2 vss vdd wl_n wl_drive
Mnmos1 vss wl_n wl_drive vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mnmos2 wl_drive wl_n vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mpmos1 vdd wl_n wl_drive vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
Mpmos2 wl_drive wl_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
.ends DP8TWLDrive_30LN100WN30LP200WP_wl2

* DP8TArray_128X32
.subckt DP8TArray_128X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
Xinst1x0 vss vdd wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
.ends DP8TArray_128X32

* DP8TArray_64X32
.subckt DP8TArray_64X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
Xinst1x0 vss vdd wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
.ends DP8TArray_64X32

* DP8TArray_32X32
.subckt DP8TArray_32X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_32X16
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X16
.ends DP8TArray_32X32

* DP8TArray_32X16
.subckt DP8TArray_32X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
Xinst1x0 vss vdd wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
.ends DP8TArray_32X16

* DP8TArray_16X16
.subckt DP8TArray_16X16 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_16X8
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X8
.ends DP8TArray_16X16

* DP8TArray_16X8
.subckt DP8TArray_16X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
.ends DP8TArray_16X8

* DP8TArray_8X8
.subckt DP8TArray_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X4
.ends DP8TArray_8X8

* DP8TArray_8X4
.subckt DP8TArray_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
.ends DP8TArray_8X4

* DP8TArray_4X4
.subckt DP8TArray_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X2
.ends DP8TArray_4X4

* DP8TArray_4X2
.subckt DP8TArray_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
.ends DP8TArray_4X2

* DP8TArray_2X2
.subckt DP8TArray_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TArray_2X1
Xinst0x1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X1
.ends DP8TArray_2X2

* DP8TArray_2X1
.subckt DP8TArray_2X1 vss vdd wl1[0] wl1[1] wl2[0] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 vdd vss wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
Xinst1x0 vdd vss wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
.ends DP8TArray_2X1

* DP8TColumnPeriphery_8B4M_bl1
.subckt DP8TColumnPeriphery_8B4M_bl1 vss vdd clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd bl[0] bl_n[0] precharge_n DP8TPrecharge_bl1
Xprecharge[1] vdd bl[1] bl_n[1] precharge_n DP8TPrecharge_bl1
Xprecharge[2] vdd bl[2] bl_n[2] precharge_n DP8TPrecharge_bl1
Xprecharge[3] vdd bl[3] bl_n[3] precharge_n DP8TPrecharge_bl1
Xprecharge[4] vdd bl[4] bl_n[4] precharge_n DP8TPrecharge_bl1
Xprecharge[5] vdd bl[5] bl_n[5] precharge_n DP8TPrecharge_bl1
Xprecharge[6] vdd bl[6] bl_n[6] precharge_n DP8TPrecharge_bl1
Xprecharge[7] vdd bl[7] bl_n[7] precharge_n DP8TPrecharge_bl1
Xprecharge[8] vdd bl[8] bl_n[8] precharge_n DP8TPrecharge_bl1
Xprecharge[9] vdd bl[9] bl_n[9] precharge_n DP8TPrecharge_bl1
Xprecharge[10] vdd bl[10] bl_n[10] precharge_n DP8TPrecharge_bl1
Xprecharge[11] vdd bl[11] bl_n[11] precharge_n DP8TPrecharge_bl1
Xprecharge[12] vdd bl[12] bl_n[12] precharge_n DP8TPrecharge_bl1
Xprecharge[13] vdd bl[13] bl_n[13] precharge_n DP8TPrecharge_bl1
Xprecharge[14] vdd bl[14] bl_n[14] precharge_n DP8TPrecharge_bl1
Xprecharge[15] vdd bl[15] bl_n[15] precharge_n DP8TPrecharge_bl1
Xprecharge[16] vdd bl[16] bl_n[16] precharge_n DP8TPrecharge_bl1
Xprecharge[17] vdd bl[17] bl_n[17] precharge_n DP8TPrecharge_bl1
Xprecharge[18] vdd bl[18] bl_n[18] precharge_n DP8TPrecharge_bl1
Xprecharge[19] vdd bl[19] bl_n[19] precharge_n DP8TPrecharge_bl1
Xprecharge[20] vdd bl[20] bl_n[20] precharge_n DP8TPrecharge_bl1
Xprecharge[21] vdd bl[21] bl_n[21] precharge_n DP8TPrecharge_bl1
Xprecharge[22] vdd bl[22] bl_n[22] precharge_n DP8TPrecharge_bl1
Xprecharge[23] vdd bl[23] bl_n[23] precharge_n DP8TPrecharge_bl1
Xprecharge[24] vdd bl[24] bl_n[24] precharge_n DP8TPrecharge_bl1
Xprecharge[25] vdd bl[25] bl_n[25] precharge_n DP8TPrecharge_bl1
Xprecharge[26] vdd bl[26] bl_n[26] precharge_n DP8TPrecharge_bl1
Xprecharge[27] vdd bl[27] bl_n[27] precharge_n DP8TPrecharge_bl1
Xprecharge[28] vdd bl[28] bl_n[28] precharge_n DP8TPrecharge_bl1
Xprecharge[29] vdd bl[29] bl_n[29] precharge_n DP8TPrecharge_bl1
Xprecharge[30] vdd bl[30] bl_n[30] precharge_n DP8TPrecharge_bl1
Xprecharge[31] vdd bl[31] bl_n[31] precharge_n DP8TPrecharge_bl1
Xcolmux[0] bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl[0] muxbl_n[0] DP8TColMux_4C_bl1
Xcolmux[1] bl[4] bl_n[4] mux[0] bl[5] bl_n[5] mux[1] bl[6] bl_n[6] mux[2] bl[7] bl_n[7] mux[3] vss muxbl[1] muxbl_n[1] DP8TColMux_4C_bl1
Xcolmux[2] bl[8] bl_n[8] mux[0] bl[9] bl_n[9] mux[1] bl[10] bl_n[10] mux[2] bl[11] bl_n[11] mux[3] vss muxbl[2] muxbl_n[2] DP8TColMux_4C_bl1
Xcolmux[3] bl[12] bl_n[12] mux[0] bl[13] bl_n[13] mux[1] bl[14] bl_n[14] mux[2] bl[15] bl_n[15] mux[3] vss muxbl[3] muxbl_n[3] DP8TColMux_4C_bl1
Xcolmux[4] bl[16] bl_n[16] mux[0] bl[17] bl_n[17] mux[1] bl[18] bl_n[18] mux[2] bl[19] bl_n[19] mux[3] vss muxbl[4] muxbl_n[4] DP8TColMux_4C_bl1
Xcolmux[5] bl[20] bl_n[20] mux[0] bl[21] bl_n[21] mux[1] bl[22] bl_n[22] mux[2] bl[23] bl_n[23] mux[3] vss muxbl[5] muxbl_n[5] DP8TColMux_4C_bl1
Xcolmux[6] bl[24] bl_n[24] mux[0] bl[25] bl_n[25] mux[1] bl[26] bl_n[26] mux[2] bl[27] bl_n[27] mux[3] vss muxbl[6] muxbl_n[6] DP8TColMux_4C_bl1
Xcolmux[7] bl[28] bl_n[28] mux[0] bl[29] bl_n[29] mux[1] bl[30] bl_n[30] mux[2] bl[31] bl_n[31] mux[3] vss muxbl[7] muxbl_n[7] DP8TColMux_4C_bl1
Xsenseamp[0] vss vdd muxbl[0] muxbl_n[0] q[0] DP8TSenseAmp_4M
Xsenseamp[1] vss vdd muxbl[1] muxbl_n[1] q[1] DP8TSenseAmp_4M
Xsenseamp[2] vss vdd muxbl[2] muxbl_n[2] q[2] DP8TSenseAmp_4M
Xsenseamp[3] vss vdd muxbl[3] muxbl_n[3] q[3] DP8TSenseAmp_4M
Xsenseamp[4] vss vdd muxbl[4] muxbl_n[4] q[4] DP8TSenseAmp_4M
Xsenseamp[5] vss vdd muxbl[5] muxbl_n[5] q[5] DP8TSenseAmp_4M
Xsenseamp[6] vss vdd muxbl[6] muxbl_n[6] q[6] DP8TSenseAmp_4M
Xsenseamp[7] vss vdd muxbl[7] muxbl_n[7] q[7] DP8TSenseAmp_4M
Xwritedrive[0] vss vdd intclk we_n muxbl[0] muxbl_n[0] d[0] muxbl[1] muxbl_n[1] d[1] DP8TWriteDriver_4M2B
Xwritedrive[1] vss vdd intclk we_n muxbl[2] muxbl_n[2] d[2] muxbl[3] muxbl_n[3] d[3] DP8TWriteDriver_4M2B
Xwritedrive[2] vss vdd intclk we_n muxbl[4] muxbl_n[4] d[4] muxbl[5] muxbl_n[5] d[5] DP8TWriteDriver_4M2B
Xwritedrive[3] vss vdd intclk we_n muxbl[6] muxbl_n[6] d[6] muxbl[7] muxbl_n[7] d[7] DP8TWriteDriver_4M2B
Xclkwe vss vdd clk intclk we we_en we_n DP8TClockWE
.ends DP8TColumnPeriphery_8B4M_bl1

* DP8TPrecharge_bl1
.subckt DP8TPrecharge_bl1 vdd bl bl_n precharge_n
Mpc1 vdd precharge_n bl vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc2 bl precharge_n bl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc3 bl_n precharge_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
.ends DP8TPrecharge_bl1

* DP8TColMux_4C_bl1
.subckt DP8TColMux_4C_bl1 bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl muxbl_n
Mpgbl0 bl[0] mux[0] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln0 muxbl_n mux[0] bl_n[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl1 bl[1] mux[1] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln1 muxbl_n mux[1] bl_n[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl2 bl[2] mux[2] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln2 muxbl_n mux[2] bl_n[2] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl3 bl[3] mux[3] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln3 muxbl_n mux[3] bl_n[3] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
.ends DP8TColMux_4C_bl1

* DP8TSenseAmp_4M
.subckt DP8TSenseAmp_4M vss vdd bl bl_n q
Xlatch vss nq q vdd bl bl_n nsnrlatch_x1
Xtie vdd vss tie
.ends DP8TSenseAmp_4M

* DP8TWriteDriver_4M2B
.subckt DP8TWriteDriver_4M2B vss vdd clk we_n bl[0] bl_n[0] d[0] bl[1] bl_n[1] d[1]
Xff[0] vdd clk vss d[0] d_latched[0] sff1_x4
Xff[1] vdd clk vss d[1] d_latched[1] sff1_x4
Xnora[0] vdd vss bl_drive[0] d_latched[0] we_n nor2_x0
Xnora[1] vdd vss bl_drive[1] d_latched[1] we_n nor2_x0
Xinv[0] vdd vss d_latched[0] d_n[0] inv_x0
Xinv[1] vdd vss d_latched[1] d_n[1] inv_x0
Xnorb[0] vdd vss bln_drive[0] d_n[0] we_n nor2_x0
Xnorb[1] vdd vss bln_drive[1] d_n[1] we_n nor2_x0
Mblpd[0] vss bl_drive[0] bl[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblpd[1] vss bl_drive[1] bl[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[0] bl_n[0] bln_drive[0] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
Mblnpd[1] bl_n[1] bln_drive[1] vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.9um
.ends DP8TWriteDriver_4M2B

* DP8TClockWE
.subckt DP8TClockWE vss vdd clkup clklow we we_en we_n
Xclkbuf vdd vss clkup clklow buf_x2
Xweff vdd clklow vss we we_latched sff1_x4
Xwenand vdd vss we_n we_en we_latched nand2_x0
.ends DP8TClockWE

* DP8TColumnPeriphery_8B4M_bl2
.subckt DP8TColumnPeriphery_8B4M_bl2 vss vdd clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd bl[0] bl_n[0] precharge_n DP8TPrecharge_bl2
Xprecharge[1] vdd bl[1] bl_n[1] precharge_n DP8TPrecharge_bl2
Xprecharge[2] vdd bl[2] bl_n[2] precharge_n DP8TPrecharge_bl2
Xprecharge[3] vdd bl[3] bl_n[3] precharge_n DP8TPrecharge_bl2
Xprecharge[4] vdd bl[4] bl_n[4] precharge_n DP8TPrecharge_bl2
Xprecharge[5] vdd bl[5] bl_n[5] precharge_n DP8TPrecharge_bl2
Xprecharge[6] vdd bl[6] bl_n[6] precharge_n DP8TPrecharge_bl2
Xprecharge[7] vdd bl[7] bl_n[7] precharge_n DP8TPrecharge_bl2
Xprecharge[8] vdd bl[8] bl_n[8] precharge_n DP8TPrecharge_bl2
Xprecharge[9] vdd bl[9] bl_n[9] precharge_n DP8TPrecharge_bl2
Xprecharge[10] vdd bl[10] bl_n[10] precharge_n DP8TPrecharge_bl2
Xprecharge[11] vdd bl[11] bl_n[11] precharge_n DP8TPrecharge_bl2
Xprecharge[12] vdd bl[12] bl_n[12] precharge_n DP8TPrecharge_bl2
Xprecharge[13] vdd bl[13] bl_n[13] precharge_n DP8TPrecharge_bl2
Xprecharge[14] vdd bl[14] bl_n[14] precharge_n DP8TPrecharge_bl2
Xprecharge[15] vdd bl[15] bl_n[15] precharge_n DP8TPrecharge_bl2
Xprecharge[16] vdd bl[16] bl_n[16] precharge_n DP8TPrecharge_bl2
Xprecharge[17] vdd bl[17] bl_n[17] precharge_n DP8TPrecharge_bl2
Xprecharge[18] vdd bl[18] bl_n[18] precharge_n DP8TPrecharge_bl2
Xprecharge[19] vdd bl[19] bl_n[19] precharge_n DP8TPrecharge_bl2
Xprecharge[20] vdd bl[20] bl_n[20] precharge_n DP8TPrecharge_bl2
Xprecharge[21] vdd bl[21] bl_n[21] precharge_n DP8TPrecharge_bl2
Xprecharge[22] vdd bl[22] bl_n[22] precharge_n DP8TPrecharge_bl2
Xprecharge[23] vdd bl[23] bl_n[23] precharge_n DP8TPrecharge_bl2
Xprecharge[24] vdd bl[24] bl_n[24] precharge_n DP8TPrecharge_bl2
Xprecharge[25] vdd bl[25] bl_n[25] precharge_n DP8TPrecharge_bl2
Xprecharge[26] vdd bl[26] bl_n[26] precharge_n DP8TPrecharge_bl2
Xprecharge[27] vdd bl[27] bl_n[27] precharge_n DP8TPrecharge_bl2
Xprecharge[28] vdd bl[28] bl_n[28] precharge_n DP8TPrecharge_bl2
Xprecharge[29] vdd bl[29] bl_n[29] precharge_n DP8TPrecharge_bl2
Xprecharge[30] vdd bl[30] bl_n[30] precharge_n DP8TPrecharge_bl2
Xprecharge[31] vdd bl[31] bl_n[31] precharge_n DP8TPrecharge_bl2
Xcolmux[0] bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl[0] muxbl_n[0] DP8TColMux_4C_bl2
Xcolmux[1] bl[4] bl_n[4] mux[0] bl[5] bl_n[5] mux[1] bl[6] bl_n[6] mux[2] bl[7] bl_n[7] mux[3] vss muxbl[1] muxbl_n[1] DP8TColMux_4C_bl2
Xcolmux[2] bl[8] bl_n[8] mux[0] bl[9] bl_n[9] mux[1] bl[10] bl_n[10] mux[2] bl[11] bl_n[11] mux[3] vss muxbl[2] muxbl_n[2] DP8TColMux_4C_bl2
Xcolmux[3] bl[12] bl_n[12] mux[0] bl[13] bl_n[13] mux[1] bl[14] bl_n[14] mux[2] bl[15] bl_n[15] mux[3] vss muxbl[3] muxbl_n[3] DP8TColMux_4C_bl2
Xcolmux[4] bl[16] bl_n[16] mux[0] bl[17] bl_n[17] mux[1] bl[18] bl_n[18] mux[2] bl[19] bl_n[19] mux[3] vss muxbl[4] muxbl_n[4] DP8TColMux_4C_bl2
Xcolmux[5] bl[20] bl_n[20] mux[0] bl[21] bl_n[21] mux[1] bl[22] bl_n[22] mux[2] bl[23] bl_n[23] mux[3] vss muxbl[5] muxbl_n[5] DP8TColMux_4C_bl2
Xcolmux[6] bl[24] bl_n[24] mux[0] bl[25] bl_n[25] mux[1] bl[26] bl_n[26] mux[2] bl[27] bl_n[27] mux[3] vss muxbl[6] muxbl_n[6] DP8TColMux_4C_bl2
Xcolmux[7] bl[28] bl_n[28] mux[0] bl[29] bl_n[29] mux[1] bl[30] bl_n[30] mux[2] bl[31] bl_n[31] mux[3] vss muxbl[7] muxbl_n[7] DP8TColMux_4C_bl2
Xsenseamp[0] vss vdd muxbl[0] muxbl_n[0] q[0] DP8TSenseAmp_4M
Xsenseamp[1] vss vdd muxbl[1] muxbl_n[1] q[1] DP8TSenseAmp_4M
Xsenseamp[2] vss vdd muxbl[2] muxbl_n[2] q[2] DP8TSenseAmp_4M
Xsenseamp[3] vss vdd muxbl[3] muxbl_n[3] q[3] DP8TSenseAmp_4M
Xsenseamp[4] vss vdd muxbl[4] muxbl_n[4] q[4] DP8TSenseAmp_4M
Xsenseamp[5] vss vdd muxbl[5] muxbl_n[5] q[5] DP8TSenseAmp_4M
Xsenseamp[6] vss vdd muxbl[6] muxbl_n[6] q[6] DP8TSenseAmp_4M
Xsenseamp[7] vss vdd muxbl[7] muxbl_n[7] q[7] DP8TSenseAmp_4M
Xwritedrive[0] vss vdd intclk we_n muxbl[0] muxbl_n[0] d[0] muxbl[1] muxbl_n[1] d[1] DP8TWriteDriver_4M2B
Xwritedrive[1] vss vdd intclk we_n muxbl[2] muxbl_n[2] d[2] muxbl[3] muxbl_n[3] d[3] DP8TWriteDriver_4M2B
Xwritedrive[2] vss vdd intclk we_n muxbl[4] muxbl_n[4] d[4] muxbl[5] muxbl_n[5] d[5] DP8TWriteDriver_4M2B
Xwritedrive[3] vss vdd intclk we_n muxbl[6] muxbl_n[6] d[6] muxbl[7] muxbl_n[7] d[7] DP8TWriteDriver_4M2B
Xclkwe vss vdd clk intclk we we_en we_n DP8TClockWE
.ends DP8TColumnPeriphery_8B4M_bl2

* DP8TPrecharge_bl2
.subckt DP8TPrecharge_bl2 vdd bl bl_n precharge_n
Mpc1 vdd precharge_n bl vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc2 bl precharge_n bl_n vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
Mpc3 bl_n precharge_n vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=0.42um
.ends DP8TPrecharge_bl2

* DP8TColMux_4C_bl2
.subckt DP8TColMux_4C_bl2 bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl muxbl_n
Mpgbl0 bl[0] mux[0] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln0 muxbl_n mux[0] bl_n[0] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl1 bl[1] mux[1] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln1 muxbl_n mux[1] bl_n[1] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl2 bl[2] mux[2] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln2 muxbl_n mux[2] bl_n[2] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbl3 bl[3] mux[3] muxbl vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
Mpgbln3 muxbl_n mux[3] bl_n[3] vss sky130_fd_pr__nfet_01v8__model l=0.15um w=4.0um
.ends DP8TColMux_4C_bl2
