-- no model for nor3_x0
