../rtl/type_dec.vhdl