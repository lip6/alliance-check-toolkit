* npn_f
.param
+ dkisnpn1x1=1.2882e+00 dkbfnpn1x1=1.5018e-00
+ dkisnpn1x2=1.3275e+00 dkbfnpn1x2=1.4758e+00
+ dkisnpnpolyhv=1.69 dkbfnpnpolyhv=1.525
