* Spice description of noa3ao322_x1
* Spice driver version -1308426469
* Date ( dd/mm/yyyy hh:mm:ss ):  2/05/2024 at 11:28:14

* INTERF i0 i1 i2 i3 i4 i5 i6 nq vdd vss 


.subckt noa3ao322_x1 13 14 9 7 6 5 8 10 4 16 
* NET 4 = vdd
* NET 5 = i5
* NET 6 = i4
* NET 7 = i3
* NET 8 = i6
* NET 9 = i2
* NET 10 = nq
* NET 13 = i0
* NET 14 = i1
* NET 16 = vss
Mtr_00014 3 5 1 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00013 1 6 2 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00012 2 7 10 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00011 10 8 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00010 3 9 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00009 4 14 3 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00008 3 13 4 4 sky130_fd_pr__pfet_01v8__model L=0.15U W=3.31U AS=0.7944P AD=0.7944P PS=7.11U PD=7.11U 
Mtr_00007 16 5 12 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00006 12 6 16 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00005 16 7 12 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00004 12 8 10 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00003 15 13 16 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00002 11 14 15 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
Mtr_00001 10 9 11 16 sky130_fd_pr__nfet_01v8__model L=0.15U W=2.04U AS=0.4896P AD=0.4896P PS=4.56U PD=4.56U 
C14 3 16 1.20336e-15
C13 4 16 2.6012e-15
C12 5 16 1.64189e-15
C11 6 16 1.70741e-15
C10 7 16 1.68002e-15
C9 8 16 1.29385e-15
C8 9 16 1.59788e-15
C7 10 16 1.85113e-15
C5 12 16 5.59015e-16
C4 13 16 1.59788e-15
C3 14 16 1.92016e-15
C1 16 16 2.8047e-15
.ends noa3ao322_x1

